module KeySchedule(
  input  [127:0] io_keyIn_bits, // @[src/main/scala/crypto/aes/KeySchedule.scala 12:14]
  output [127:0] io_rks_0_bits, // @[src/main/scala/crypto/aes/KeySchedule.scala 12:14]
  output [127:0] io_rks_1_bits, // @[src/main/scala/crypto/aes/KeySchedule.scala 12:14]
  output [127:0] io_rks_2_bits, // @[src/main/scala/crypto/aes/KeySchedule.scala 12:14]
  output [127:0] io_rks_3_bits, // @[src/main/scala/crypto/aes/KeySchedule.scala 12:14]
  output [127:0] io_rks_4_bits, // @[src/main/scala/crypto/aes/KeySchedule.scala 12:14]
  output [127:0] io_rks_5_bits, // @[src/main/scala/crypto/aes/KeySchedule.scala 12:14]
  output [127:0] io_rks_6_bits, // @[src/main/scala/crypto/aes/KeySchedule.scala 12:14]
  output [127:0] io_rks_7_bits, // @[src/main/scala/crypto/aes/KeySchedule.scala 12:14]
  output [127:0] io_rks_8_bits, // @[src/main/scala/crypto/aes/KeySchedule.scala 12:14]
  output [127:0] io_rks_9_bits, // @[src/main/scala/crypto/aes/KeySchedule.scala 12:14]
  output [127:0] io_rks_10_bits // @[src/main/scala/crypto/aes/KeySchedule.scala 12:14]
);
  wire [31:0] w_0 = io_keyIn_bits[127:96]; // @[src/main/scala/crypto/aes/KeySchedule.scala 49:26]
  wire [31:0] w_1 = io_keyIn_bits[95:64]; // @[src/main/scala/crypto/aes/KeySchedule.scala 49:26]
  wire [31:0] w_2 = io_keyIn_bits[63:32]; // @[src/main/scala/crypto/aes/KeySchedule.scala 49:26]
  wire [31:0] w_3 = io_keyIn_bits[31:0]; // @[src/main/scala/crypto/aes/KeySchedule.scala 49:26]
  wire [31:0] _t_T_2 = {w_3[23:0],w_3[31:24]}; // @[src/main/scala/crypto/aes/KeySchedule.scala 23:43]
  wire [7:0] _GEN_1 = 8'h1 == _t_T_2[15:8] ? 8'h7c : 8'h63; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2 = 8'h2 == _t_T_2[15:8] ? 8'h77 : _GEN_1; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3 = 8'h3 == _t_T_2[15:8] ? 8'h7b : _GEN_2; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4 = 8'h4 == _t_T_2[15:8] ? 8'hf2 : _GEN_3; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5 = 8'h5 == _t_T_2[15:8] ? 8'h6b : _GEN_4; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6 = 8'h6 == _t_T_2[15:8] ? 8'h6f : _GEN_5; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7 = 8'h7 == _t_T_2[15:8] ? 8'hc5 : _GEN_6; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8 = 8'h8 == _t_T_2[15:8] ? 8'h30 : _GEN_7; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9 = 8'h9 == _t_T_2[15:8] ? 8'h1 : _GEN_8; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10 = 8'ha == _t_T_2[15:8] ? 8'h67 : _GEN_9; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_11 = 8'hb == _t_T_2[15:8] ? 8'h2b : _GEN_10; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_12 = 8'hc == _t_T_2[15:8] ? 8'hfe : _GEN_11; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_13 = 8'hd == _t_T_2[15:8] ? 8'hd7 : _GEN_12; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_14 = 8'he == _t_T_2[15:8] ? 8'hab : _GEN_13; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_15 = 8'hf == _t_T_2[15:8] ? 8'h76 : _GEN_14; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_16 = 8'h10 == _t_T_2[15:8] ? 8'hca : _GEN_15; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_17 = 8'h11 == _t_T_2[15:8] ? 8'h82 : _GEN_16; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_18 = 8'h12 == _t_T_2[15:8] ? 8'hc9 : _GEN_17; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_19 = 8'h13 == _t_T_2[15:8] ? 8'h7d : _GEN_18; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_20 = 8'h14 == _t_T_2[15:8] ? 8'hfa : _GEN_19; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_21 = 8'h15 == _t_T_2[15:8] ? 8'h59 : _GEN_20; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_22 = 8'h16 == _t_T_2[15:8] ? 8'h47 : _GEN_21; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_23 = 8'h17 == _t_T_2[15:8] ? 8'hf0 : _GEN_22; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_24 = 8'h18 == _t_T_2[15:8] ? 8'had : _GEN_23; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_25 = 8'h19 == _t_T_2[15:8] ? 8'hd4 : _GEN_24; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_26 = 8'h1a == _t_T_2[15:8] ? 8'ha2 : _GEN_25; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_27 = 8'h1b == _t_T_2[15:8] ? 8'haf : _GEN_26; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_28 = 8'h1c == _t_T_2[15:8] ? 8'h9c : _GEN_27; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_29 = 8'h1d == _t_T_2[15:8] ? 8'ha4 : _GEN_28; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_30 = 8'h1e == _t_T_2[15:8] ? 8'h72 : _GEN_29; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_31 = 8'h1f == _t_T_2[15:8] ? 8'hc0 : _GEN_30; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_32 = 8'h20 == _t_T_2[15:8] ? 8'hb7 : _GEN_31; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_33 = 8'h21 == _t_T_2[15:8] ? 8'hfd : _GEN_32; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_34 = 8'h22 == _t_T_2[15:8] ? 8'h93 : _GEN_33; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_35 = 8'h23 == _t_T_2[15:8] ? 8'h26 : _GEN_34; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_36 = 8'h24 == _t_T_2[15:8] ? 8'h36 : _GEN_35; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_37 = 8'h25 == _t_T_2[15:8] ? 8'h3f : _GEN_36; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_38 = 8'h26 == _t_T_2[15:8] ? 8'hf7 : _GEN_37; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_39 = 8'h27 == _t_T_2[15:8] ? 8'hcc : _GEN_38; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_40 = 8'h28 == _t_T_2[15:8] ? 8'h34 : _GEN_39; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_41 = 8'h29 == _t_T_2[15:8] ? 8'ha5 : _GEN_40; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_42 = 8'h2a == _t_T_2[15:8] ? 8'he5 : _GEN_41; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_43 = 8'h2b == _t_T_2[15:8] ? 8'hf1 : _GEN_42; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_44 = 8'h2c == _t_T_2[15:8] ? 8'h71 : _GEN_43; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_45 = 8'h2d == _t_T_2[15:8] ? 8'hd8 : _GEN_44; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_46 = 8'h2e == _t_T_2[15:8] ? 8'h31 : _GEN_45; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_47 = 8'h2f == _t_T_2[15:8] ? 8'h15 : _GEN_46; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_48 = 8'h30 == _t_T_2[15:8] ? 8'h4 : _GEN_47; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_49 = 8'h31 == _t_T_2[15:8] ? 8'hc7 : _GEN_48; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_50 = 8'h32 == _t_T_2[15:8] ? 8'h23 : _GEN_49; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_51 = 8'h33 == _t_T_2[15:8] ? 8'hc3 : _GEN_50; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_52 = 8'h34 == _t_T_2[15:8] ? 8'h18 : _GEN_51; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_53 = 8'h35 == _t_T_2[15:8] ? 8'h96 : _GEN_52; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_54 = 8'h36 == _t_T_2[15:8] ? 8'h5 : _GEN_53; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_55 = 8'h37 == _t_T_2[15:8] ? 8'h9a : _GEN_54; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_56 = 8'h38 == _t_T_2[15:8] ? 8'h7 : _GEN_55; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_57 = 8'h39 == _t_T_2[15:8] ? 8'h12 : _GEN_56; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_58 = 8'h3a == _t_T_2[15:8] ? 8'h80 : _GEN_57; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_59 = 8'h3b == _t_T_2[15:8] ? 8'he2 : _GEN_58; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_60 = 8'h3c == _t_T_2[15:8] ? 8'heb : _GEN_59; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_61 = 8'h3d == _t_T_2[15:8] ? 8'h27 : _GEN_60; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_62 = 8'h3e == _t_T_2[15:8] ? 8'hb2 : _GEN_61; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_63 = 8'h3f == _t_T_2[15:8] ? 8'h75 : _GEN_62; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_64 = 8'h40 == _t_T_2[15:8] ? 8'h9 : _GEN_63; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_65 = 8'h41 == _t_T_2[15:8] ? 8'h83 : _GEN_64; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_66 = 8'h42 == _t_T_2[15:8] ? 8'h2c : _GEN_65; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_67 = 8'h43 == _t_T_2[15:8] ? 8'h1a : _GEN_66; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_68 = 8'h44 == _t_T_2[15:8] ? 8'h1b : _GEN_67; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_69 = 8'h45 == _t_T_2[15:8] ? 8'h6e : _GEN_68; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_70 = 8'h46 == _t_T_2[15:8] ? 8'h5a : _GEN_69; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_71 = 8'h47 == _t_T_2[15:8] ? 8'ha0 : _GEN_70; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_72 = 8'h48 == _t_T_2[15:8] ? 8'h52 : _GEN_71; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_73 = 8'h49 == _t_T_2[15:8] ? 8'h3b : _GEN_72; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_74 = 8'h4a == _t_T_2[15:8] ? 8'hd6 : _GEN_73; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_75 = 8'h4b == _t_T_2[15:8] ? 8'hb3 : _GEN_74; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_76 = 8'h4c == _t_T_2[15:8] ? 8'h29 : _GEN_75; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_77 = 8'h4d == _t_T_2[15:8] ? 8'he3 : _GEN_76; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_78 = 8'h4e == _t_T_2[15:8] ? 8'h2f : _GEN_77; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_79 = 8'h4f == _t_T_2[15:8] ? 8'h84 : _GEN_78; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_80 = 8'h50 == _t_T_2[15:8] ? 8'h53 : _GEN_79; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_81 = 8'h51 == _t_T_2[15:8] ? 8'hd1 : _GEN_80; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_82 = 8'h52 == _t_T_2[15:8] ? 8'h0 : _GEN_81; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_83 = 8'h53 == _t_T_2[15:8] ? 8'hed : _GEN_82; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_84 = 8'h54 == _t_T_2[15:8] ? 8'h20 : _GEN_83; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_85 = 8'h55 == _t_T_2[15:8] ? 8'hfc : _GEN_84; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_86 = 8'h56 == _t_T_2[15:8] ? 8'hb1 : _GEN_85; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_87 = 8'h57 == _t_T_2[15:8] ? 8'h5b : _GEN_86; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_88 = 8'h58 == _t_T_2[15:8] ? 8'h6a : _GEN_87; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_89 = 8'h59 == _t_T_2[15:8] ? 8'hcb : _GEN_88; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_90 = 8'h5a == _t_T_2[15:8] ? 8'hbe : _GEN_89; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_91 = 8'h5b == _t_T_2[15:8] ? 8'h39 : _GEN_90; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_92 = 8'h5c == _t_T_2[15:8] ? 8'h4a : _GEN_91; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_93 = 8'h5d == _t_T_2[15:8] ? 8'h4c : _GEN_92; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_94 = 8'h5e == _t_T_2[15:8] ? 8'h58 : _GEN_93; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_95 = 8'h5f == _t_T_2[15:8] ? 8'hcf : _GEN_94; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_96 = 8'h60 == _t_T_2[15:8] ? 8'hd0 : _GEN_95; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_97 = 8'h61 == _t_T_2[15:8] ? 8'hef : _GEN_96; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_98 = 8'h62 == _t_T_2[15:8] ? 8'haa : _GEN_97; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_99 = 8'h63 == _t_T_2[15:8] ? 8'hfb : _GEN_98; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_100 = 8'h64 == _t_T_2[15:8] ? 8'h43 : _GEN_99; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_101 = 8'h65 == _t_T_2[15:8] ? 8'h4d : _GEN_100; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_102 = 8'h66 == _t_T_2[15:8] ? 8'h33 : _GEN_101; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_103 = 8'h67 == _t_T_2[15:8] ? 8'h85 : _GEN_102; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_104 = 8'h68 == _t_T_2[15:8] ? 8'h45 : _GEN_103; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_105 = 8'h69 == _t_T_2[15:8] ? 8'hf9 : _GEN_104; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_106 = 8'h6a == _t_T_2[15:8] ? 8'h2 : _GEN_105; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_107 = 8'h6b == _t_T_2[15:8] ? 8'h7f : _GEN_106; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_108 = 8'h6c == _t_T_2[15:8] ? 8'h50 : _GEN_107; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_109 = 8'h6d == _t_T_2[15:8] ? 8'h3c : _GEN_108; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_110 = 8'h6e == _t_T_2[15:8] ? 8'h9f : _GEN_109; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_111 = 8'h6f == _t_T_2[15:8] ? 8'ha8 : _GEN_110; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_112 = 8'h70 == _t_T_2[15:8] ? 8'h51 : _GEN_111; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_113 = 8'h71 == _t_T_2[15:8] ? 8'ha3 : _GEN_112; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_114 = 8'h72 == _t_T_2[15:8] ? 8'h40 : _GEN_113; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_115 = 8'h73 == _t_T_2[15:8] ? 8'h8f : _GEN_114; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_116 = 8'h74 == _t_T_2[15:8] ? 8'h92 : _GEN_115; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_117 = 8'h75 == _t_T_2[15:8] ? 8'h9d : _GEN_116; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_118 = 8'h76 == _t_T_2[15:8] ? 8'h38 : _GEN_117; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_119 = 8'h77 == _t_T_2[15:8] ? 8'hf5 : _GEN_118; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_120 = 8'h78 == _t_T_2[15:8] ? 8'hbc : _GEN_119; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_121 = 8'h79 == _t_T_2[15:8] ? 8'hb6 : _GEN_120; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_122 = 8'h7a == _t_T_2[15:8] ? 8'hda : _GEN_121; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_123 = 8'h7b == _t_T_2[15:8] ? 8'h21 : _GEN_122; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_124 = 8'h7c == _t_T_2[15:8] ? 8'h10 : _GEN_123; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_125 = 8'h7d == _t_T_2[15:8] ? 8'hff : _GEN_124; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_126 = 8'h7e == _t_T_2[15:8] ? 8'hf3 : _GEN_125; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_127 = 8'h7f == _t_T_2[15:8] ? 8'hd2 : _GEN_126; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_128 = 8'h80 == _t_T_2[15:8] ? 8'hcd : _GEN_127; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_129 = 8'h81 == _t_T_2[15:8] ? 8'hc : _GEN_128; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_130 = 8'h82 == _t_T_2[15:8] ? 8'h13 : _GEN_129; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_131 = 8'h83 == _t_T_2[15:8] ? 8'hec : _GEN_130; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_132 = 8'h84 == _t_T_2[15:8] ? 8'h5f : _GEN_131; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_133 = 8'h85 == _t_T_2[15:8] ? 8'h97 : _GEN_132; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_134 = 8'h86 == _t_T_2[15:8] ? 8'h44 : _GEN_133; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_135 = 8'h87 == _t_T_2[15:8] ? 8'h17 : _GEN_134; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_136 = 8'h88 == _t_T_2[15:8] ? 8'hc4 : _GEN_135; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_137 = 8'h89 == _t_T_2[15:8] ? 8'ha7 : _GEN_136; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_138 = 8'h8a == _t_T_2[15:8] ? 8'h7e : _GEN_137; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_139 = 8'h8b == _t_T_2[15:8] ? 8'h3d : _GEN_138; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_140 = 8'h8c == _t_T_2[15:8] ? 8'h64 : _GEN_139; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_141 = 8'h8d == _t_T_2[15:8] ? 8'h5d : _GEN_140; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_142 = 8'h8e == _t_T_2[15:8] ? 8'h19 : _GEN_141; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_143 = 8'h8f == _t_T_2[15:8] ? 8'h73 : _GEN_142; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_144 = 8'h90 == _t_T_2[15:8] ? 8'h60 : _GEN_143; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_145 = 8'h91 == _t_T_2[15:8] ? 8'h81 : _GEN_144; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_146 = 8'h92 == _t_T_2[15:8] ? 8'h4f : _GEN_145; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_147 = 8'h93 == _t_T_2[15:8] ? 8'hdc : _GEN_146; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_148 = 8'h94 == _t_T_2[15:8] ? 8'h22 : _GEN_147; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_149 = 8'h95 == _t_T_2[15:8] ? 8'h2a : _GEN_148; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_150 = 8'h96 == _t_T_2[15:8] ? 8'h90 : _GEN_149; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_151 = 8'h97 == _t_T_2[15:8] ? 8'h88 : _GEN_150; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_152 = 8'h98 == _t_T_2[15:8] ? 8'h46 : _GEN_151; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_153 = 8'h99 == _t_T_2[15:8] ? 8'hee : _GEN_152; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_154 = 8'h9a == _t_T_2[15:8] ? 8'hb8 : _GEN_153; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_155 = 8'h9b == _t_T_2[15:8] ? 8'h14 : _GEN_154; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_156 = 8'h9c == _t_T_2[15:8] ? 8'hde : _GEN_155; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_157 = 8'h9d == _t_T_2[15:8] ? 8'h5e : _GEN_156; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_158 = 8'h9e == _t_T_2[15:8] ? 8'hb : _GEN_157; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_159 = 8'h9f == _t_T_2[15:8] ? 8'hdb : _GEN_158; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_160 = 8'ha0 == _t_T_2[15:8] ? 8'he0 : _GEN_159; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_161 = 8'ha1 == _t_T_2[15:8] ? 8'h32 : _GEN_160; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_162 = 8'ha2 == _t_T_2[15:8] ? 8'h3a : _GEN_161; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_163 = 8'ha3 == _t_T_2[15:8] ? 8'ha : _GEN_162; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_164 = 8'ha4 == _t_T_2[15:8] ? 8'h49 : _GEN_163; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_165 = 8'ha5 == _t_T_2[15:8] ? 8'h6 : _GEN_164; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_166 = 8'ha6 == _t_T_2[15:8] ? 8'h24 : _GEN_165; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_167 = 8'ha7 == _t_T_2[15:8] ? 8'h5c : _GEN_166; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_168 = 8'ha8 == _t_T_2[15:8] ? 8'hc2 : _GEN_167; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_169 = 8'ha9 == _t_T_2[15:8] ? 8'hd3 : _GEN_168; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_170 = 8'haa == _t_T_2[15:8] ? 8'hac : _GEN_169; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_171 = 8'hab == _t_T_2[15:8] ? 8'h62 : _GEN_170; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_172 = 8'hac == _t_T_2[15:8] ? 8'h91 : _GEN_171; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_173 = 8'had == _t_T_2[15:8] ? 8'h95 : _GEN_172; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_174 = 8'hae == _t_T_2[15:8] ? 8'he4 : _GEN_173; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_175 = 8'haf == _t_T_2[15:8] ? 8'h79 : _GEN_174; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_176 = 8'hb0 == _t_T_2[15:8] ? 8'he7 : _GEN_175; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_177 = 8'hb1 == _t_T_2[15:8] ? 8'hc8 : _GEN_176; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_178 = 8'hb2 == _t_T_2[15:8] ? 8'h37 : _GEN_177; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_179 = 8'hb3 == _t_T_2[15:8] ? 8'h6d : _GEN_178; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_180 = 8'hb4 == _t_T_2[15:8] ? 8'h8d : _GEN_179; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_181 = 8'hb5 == _t_T_2[15:8] ? 8'hd5 : _GEN_180; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_182 = 8'hb6 == _t_T_2[15:8] ? 8'h4e : _GEN_181; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_183 = 8'hb7 == _t_T_2[15:8] ? 8'ha9 : _GEN_182; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_184 = 8'hb8 == _t_T_2[15:8] ? 8'h6c : _GEN_183; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_185 = 8'hb9 == _t_T_2[15:8] ? 8'h56 : _GEN_184; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_186 = 8'hba == _t_T_2[15:8] ? 8'hf4 : _GEN_185; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_187 = 8'hbb == _t_T_2[15:8] ? 8'hea : _GEN_186; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_188 = 8'hbc == _t_T_2[15:8] ? 8'h65 : _GEN_187; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_189 = 8'hbd == _t_T_2[15:8] ? 8'h7a : _GEN_188; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_190 = 8'hbe == _t_T_2[15:8] ? 8'hae : _GEN_189; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_191 = 8'hbf == _t_T_2[15:8] ? 8'h8 : _GEN_190; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_192 = 8'hc0 == _t_T_2[15:8] ? 8'hba : _GEN_191; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_193 = 8'hc1 == _t_T_2[15:8] ? 8'h78 : _GEN_192; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_194 = 8'hc2 == _t_T_2[15:8] ? 8'h25 : _GEN_193; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_195 = 8'hc3 == _t_T_2[15:8] ? 8'h2e : _GEN_194; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_196 = 8'hc4 == _t_T_2[15:8] ? 8'h1c : _GEN_195; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_197 = 8'hc5 == _t_T_2[15:8] ? 8'ha6 : _GEN_196; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_198 = 8'hc6 == _t_T_2[15:8] ? 8'hb4 : _GEN_197; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_199 = 8'hc7 == _t_T_2[15:8] ? 8'hc6 : _GEN_198; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_200 = 8'hc8 == _t_T_2[15:8] ? 8'he8 : _GEN_199; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_201 = 8'hc9 == _t_T_2[15:8] ? 8'hdd : _GEN_200; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_202 = 8'hca == _t_T_2[15:8] ? 8'h74 : _GEN_201; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_203 = 8'hcb == _t_T_2[15:8] ? 8'h1f : _GEN_202; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_204 = 8'hcc == _t_T_2[15:8] ? 8'h4b : _GEN_203; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_205 = 8'hcd == _t_T_2[15:8] ? 8'hbd : _GEN_204; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_206 = 8'hce == _t_T_2[15:8] ? 8'h8b : _GEN_205; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_207 = 8'hcf == _t_T_2[15:8] ? 8'h8a : _GEN_206; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_208 = 8'hd0 == _t_T_2[15:8] ? 8'h70 : _GEN_207; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_209 = 8'hd1 == _t_T_2[15:8] ? 8'h3e : _GEN_208; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_210 = 8'hd2 == _t_T_2[15:8] ? 8'hb5 : _GEN_209; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_211 = 8'hd3 == _t_T_2[15:8] ? 8'h66 : _GEN_210; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_212 = 8'hd4 == _t_T_2[15:8] ? 8'h48 : _GEN_211; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_213 = 8'hd5 == _t_T_2[15:8] ? 8'h3 : _GEN_212; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_214 = 8'hd6 == _t_T_2[15:8] ? 8'hf6 : _GEN_213; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_215 = 8'hd7 == _t_T_2[15:8] ? 8'he : _GEN_214; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_216 = 8'hd8 == _t_T_2[15:8] ? 8'h61 : _GEN_215; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_217 = 8'hd9 == _t_T_2[15:8] ? 8'h35 : _GEN_216; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_218 = 8'hda == _t_T_2[15:8] ? 8'h57 : _GEN_217; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_219 = 8'hdb == _t_T_2[15:8] ? 8'hb9 : _GEN_218; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_220 = 8'hdc == _t_T_2[15:8] ? 8'h86 : _GEN_219; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_221 = 8'hdd == _t_T_2[15:8] ? 8'hc1 : _GEN_220; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_222 = 8'hde == _t_T_2[15:8] ? 8'h1d : _GEN_221; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_223 = 8'hdf == _t_T_2[15:8] ? 8'h9e : _GEN_222; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_224 = 8'he0 == _t_T_2[15:8] ? 8'he1 : _GEN_223; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_225 = 8'he1 == _t_T_2[15:8] ? 8'hf8 : _GEN_224; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_226 = 8'he2 == _t_T_2[15:8] ? 8'h98 : _GEN_225; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_227 = 8'he3 == _t_T_2[15:8] ? 8'h11 : _GEN_226; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_228 = 8'he4 == _t_T_2[15:8] ? 8'h69 : _GEN_227; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_229 = 8'he5 == _t_T_2[15:8] ? 8'hd9 : _GEN_228; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_230 = 8'he6 == _t_T_2[15:8] ? 8'h8e : _GEN_229; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_231 = 8'he7 == _t_T_2[15:8] ? 8'h94 : _GEN_230; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_232 = 8'he8 == _t_T_2[15:8] ? 8'h9b : _GEN_231; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_233 = 8'he9 == _t_T_2[15:8] ? 8'h1e : _GEN_232; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_234 = 8'hea == _t_T_2[15:8] ? 8'h87 : _GEN_233; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_235 = 8'heb == _t_T_2[15:8] ? 8'he9 : _GEN_234; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_236 = 8'hec == _t_T_2[15:8] ? 8'hce : _GEN_235; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_237 = 8'hed == _t_T_2[15:8] ? 8'h55 : _GEN_236; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_238 = 8'hee == _t_T_2[15:8] ? 8'h28 : _GEN_237; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_239 = 8'hef == _t_T_2[15:8] ? 8'hdf : _GEN_238; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_240 = 8'hf0 == _t_T_2[15:8] ? 8'h8c : _GEN_239; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_241 = 8'hf1 == _t_T_2[15:8] ? 8'ha1 : _GEN_240; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_242 = 8'hf2 == _t_T_2[15:8] ? 8'h89 : _GEN_241; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_243 = 8'hf3 == _t_T_2[15:8] ? 8'hd : _GEN_242; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_244 = 8'hf4 == _t_T_2[15:8] ? 8'hbf : _GEN_243; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_245 = 8'hf5 == _t_T_2[15:8] ? 8'he6 : _GEN_244; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_246 = 8'hf6 == _t_T_2[15:8] ? 8'h42 : _GEN_245; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_247 = 8'hf7 == _t_T_2[15:8] ? 8'h68 : _GEN_246; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_248 = 8'hf8 == _t_T_2[15:8] ? 8'h41 : _GEN_247; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_249 = 8'hf9 == _t_T_2[15:8] ? 8'h99 : _GEN_248; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_250 = 8'hfa == _t_T_2[15:8] ? 8'h2d : _GEN_249; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_251 = 8'hfb == _t_T_2[15:8] ? 8'hf : _GEN_250; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_252 = 8'hfc == _t_T_2[15:8] ? 8'hb0 : _GEN_251; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_253 = 8'hfd == _t_T_2[15:8] ? 8'h54 : _GEN_252; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_254 = 8'hfe == _t_T_2[15:8] ? 8'hbb : _GEN_253; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_255 = 8'hff == _t_T_2[15:8] ? 8'h16 : _GEN_254; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_257 = 8'h1 == _t_T_2[7:0] ? 8'h7c : 8'h63; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_258 = 8'h2 == _t_T_2[7:0] ? 8'h77 : _GEN_257; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_259 = 8'h3 == _t_T_2[7:0] ? 8'h7b : _GEN_258; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_260 = 8'h4 == _t_T_2[7:0] ? 8'hf2 : _GEN_259; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_261 = 8'h5 == _t_T_2[7:0] ? 8'h6b : _GEN_260; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_262 = 8'h6 == _t_T_2[7:0] ? 8'h6f : _GEN_261; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_263 = 8'h7 == _t_T_2[7:0] ? 8'hc5 : _GEN_262; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_264 = 8'h8 == _t_T_2[7:0] ? 8'h30 : _GEN_263; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_265 = 8'h9 == _t_T_2[7:0] ? 8'h1 : _GEN_264; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_266 = 8'ha == _t_T_2[7:0] ? 8'h67 : _GEN_265; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_267 = 8'hb == _t_T_2[7:0] ? 8'h2b : _GEN_266; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_268 = 8'hc == _t_T_2[7:0] ? 8'hfe : _GEN_267; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_269 = 8'hd == _t_T_2[7:0] ? 8'hd7 : _GEN_268; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_270 = 8'he == _t_T_2[7:0] ? 8'hab : _GEN_269; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_271 = 8'hf == _t_T_2[7:0] ? 8'h76 : _GEN_270; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_272 = 8'h10 == _t_T_2[7:0] ? 8'hca : _GEN_271; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_273 = 8'h11 == _t_T_2[7:0] ? 8'h82 : _GEN_272; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_274 = 8'h12 == _t_T_2[7:0] ? 8'hc9 : _GEN_273; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_275 = 8'h13 == _t_T_2[7:0] ? 8'h7d : _GEN_274; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_276 = 8'h14 == _t_T_2[7:0] ? 8'hfa : _GEN_275; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_277 = 8'h15 == _t_T_2[7:0] ? 8'h59 : _GEN_276; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_278 = 8'h16 == _t_T_2[7:0] ? 8'h47 : _GEN_277; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_279 = 8'h17 == _t_T_2[7:0] ? 8'hf0 : _GEN_278; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_280 = 8'h18 == _t_T_2[7:0] ? 8'had : _GEN_279; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_281 = 8'h19 == _t_T_2[7:0] ? 8'hd4 : _GEN_280; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_282 = 8'h1a == _t_T_2[7:0] ? 8'ha2 : _GEN_281; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_283 = 8'h1b == _t_T_2[7:0] ? 8'haf : _GEN_282; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_284 = 8'h1c == _t_T_2[7:0] ? 8'h9c : _GEN_283; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_285 = 8'h1d == _t_T_2[7:0] ? 8'ha4 : _GEN_284; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_286 = 8'h1e == _t_T_2[7:0] ? 8'h72 : _GEN_285; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_287 = 8'h1f == _t_T_2[7:0] ? 8'hc0 : _GEN_286; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_288 = 8'h20 == _t_T_2[7:0] ? 8'hb7 : _GEN_287; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_289 = 8'h21 == _t_T_2[7:0] ? 8'hfd : _GEN_288; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_290 = 8'h22 == _t_T_2[7:0] ? 8'h93 : _GEN_289; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_291 = 8'h23 == _t_T_2[7:0] ? 8'h26 : _GEN_290; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_292 = 8'h24 == _t_T_2[7:0] ? 8'h36 : _GEN_291; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_293 = 8'h25 == _t_T_2[7:0] ? 8'h3f : _GEN_292; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_294 = 8'h26 == _t_T_2[7:0] ? 8'hf7 : _GEN_293; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_295 = 8'h27 == _t_T_2[7:0] ? 8'hcc : _GEN_294; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_296 = 8'h28 == _t_T_2[7:0] ? 8'h34 : _GEN_295; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_297 = 8'h29 == _t_T_2[7:0] ? 8'ha5 : _GEN_296; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_298 = 8'h2a == _t_T_2[7:0] ? 8'he5 : _GEN_297; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_299 = 8'h2b == _t_T_2[7:0] ? 8'hf1 : _GEN_298; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_300 = 8'h2c == _t_T_2[7:0] ? 8'h71 : _GEN_299; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_301 = 8'h2d == _t_T_2[7:0] ? 8'hd8 : _GEN_300; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_302 = 8'h2e == _t_T_2[7:0] ? 8'h31 : _GEN_301; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_303 = 8'h2f == _t_T_2[7:0] ? 8'h15 : _GEN_302; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_304 = 8'h30 == _t_T_2[7:0] ? 8'h4 : _GEN_303; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_305 = 8'h31 == _t_T_2[7:0] ? 8'hc7 : _GEN_304; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_306 = 8'h32 == _t_T_2[7:0] ? 8'h23 : _GEN_305; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_307 = 8'h33 == _t_T_2[7:0] ? 8'hc3 : _GEN_306; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_308 = 8'h34 == _t_T_2[7:0] ? 8'h18 : _GEN_307; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_309 = 8'h35 == _t_T_2[7:0] ? 8'h96 : _GEN_308; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_310 = 8'h36 == _t_T_2[7:0] ? 8'h5 : _GEN_309; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_311 = 8'h37 == _t_T_2[7:0] ? 8'h9a : _GEN_310; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_312 = 8'h38 == _t_T_2[7:0] ? 8'h7 : _GEN_311; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_313 = 8'h39 == _t_T_2[7:0] ? 8'h12 : _GEN_312; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_314 = 8'h3a == _t_T_2[7:0] ? 8'h80 : _GEN_313; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_315 = 8'h3b == _t_T_2[7:0] ? 8'he2 : _GEN_314; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_316 = 8'h3c == _t_T_2[7:0] ? 8'heb : _GEN_315; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_317 = 8'h3d == _t_T_2[7:0] ? 8'h27 : _GEN_316; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_318 = 8'h3e == _t_T_2[7:0] ? 8'hb2 : _GEN_317; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_319 = 8'h3f == _t_T_2[7:0] ? 8'h75 : _GEN_318; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_320 = 8'h40 == _t_T_2[7:0] ? 8'h9 : _GEN_319; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_321 = 8'h41 == _t_T_2[7:0] ? 8'h83 : _GEN_320; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_322 = 8'h42 == _t_T_2[7:0] ? 8'h2c : _GEN_321; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_323 = 8'h43 == _t_T_2[7:0] ? 8'h1a : _GEN_322; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_324 = 8'h44 == _t_T_2[7:0] ? 8'h1b : _GEN_323; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_325 = 8'h45 == _t_T_2[7:0] ? 8'h6e : _GEN_324; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_326 = 8'h46 == _t_T_2[7:0] ? 8'h5a : _GEN_325; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_327 = 8'h47 == _t_T_2[7:0] ? 8'ha0 : _GEN_326; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_328 = 8'h48 == _t_T_2[7:0] ? 8'h52 : _GEN_327; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_329 = 8'h49 == _t_T_2[7:0] ? 8'h3b : _GEN_328; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_330 = 8'h4a == _t_T_2[7:0] ? 8'hd6 : _GEN_329; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_331 = 8'h4b == _t_T_2[7:0] ? 8'hb3 : _GEN_330; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_332 = 8'h4c == _t_T_2[7:0] ? 8'h29 : _GEN_331; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_333 = 8'h4d == _t_T_2[7:0] ? 8'he3 : _GEN_332; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_334 = 8'h4e == _t_T_2[7:0] ? 8'h2f : _GEN_333; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_335 = 8'h4f == _t_T_2[7:0] ? 8'h84 : _GEN_334; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_336 = 8'h50 == _t_T_2[7:0] ? 8'h53 : _GEN_335; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_337 = 8'h51 == _t_T_2[7:0] ? 8'hd1 : _GEN_336; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_338 = 8'h52 == _t_T_2[7:0] ? 8'h0 : _GEN_337; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_339 = 8'h53 == _t_T_2[7:0] ? 8'hed : _GEN_338; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_340 = 8'h54 == _t_T_2[7:0] ? 8'h20 : _GEN_339; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_341 = 8'h55 == _t_T_2[7:0] ? 8'hfc : _GEN_340; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_342 = 8'h56 == _t_T_2[7:0] ? 8'hb1 : _GEN_341; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_343 = 8'h57 == _t_T_2[7:0] ? 8'h5b : _GEN_342; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_344 = 8'h58 == _t_T_2[7:0] ? 8'h6a : _GEN_343; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_345 = 8'h59 == _t_T_2[7:0] ? 8'hcb : _GEN_344; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_346 = 8'h5a == _t_T_2[7:0] ? 8'hbe : _GEN_345; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_347 = 8'h5b == _t_T_2[7:0] ? 8'h39 : _GEN_346; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_348 = 8'h5c == _t_T_2[7:0] ? 8'h4a : _GEN_347; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_349 = 8'h5d == _t_T_2[7:0] ? 8'h4c : _GEN_348; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_350 = 8'h5e == _t_T_2[7:0] ? 8'h58 : _GEN_349; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_351 = 8'h5f == _t_T_2[7:0] ? 8'hcf : _GEN_350; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_352 = 8'h60 == _t_T_2[7:0] ? 8'hd0 : _GEN_351; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_353 = 8'h61 == _t_T_2[7:0] ? 8'hef : _GEN_352; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_354 = 8'h62 == _t_T_2[7:0] ? 8'haa : _GEN_353; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_355 = 8'h63 == _t_T_2[7:0] ? 8'hfb : _GEN_354; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_356 = 8'h64 == _t_T_2[7:0] ? 8'h43 : _GEN_355; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_357 = 8'h65 == _t_T_2[7:0] ? 8'h4d : _GEN_356; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_358 = 8'h66 == _t_T_2[7:0] ? 8'h33 : _GEN_357; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_359 = 8'h67 == _t_T_2[7:0] ? 8'h85 : _GEN_358; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_360 = 8'h68 == _t_T_2[7:0] ? 8'h45 : _GEN_359; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_361 = 8'h69 == _t_T_2[7:0] ? 8'hf9 : _GEN_360; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_362 = 8'h6a == _t_T_2[7:0] ? 8'h2 : _GEN_361; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_363 = 8'h6b == _t_T_2[7:0] ? 8'h7f : _GEN_362; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_364 = 8'h6c == _t_T_2[7:0] ? 8'h50 : _GEN_363; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_365 = 8'h6d == _t_T_2[7:0] ? 8'h3c : _GEN_364; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_366 = 8'h6e == _t_T_2[7:0] ? 8'h9f : _GEN_365; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_367 = 8'h6f == _t_T_2[7:0] ? 8'ha8 : _GEN_366; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_368 = 8'h70 == _t_T_2[7:0] ? 8'h51 : _GEN_367; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_369 = 8'h71 == _t_T_2[7:0] ? 8'ha3 : _GEN_368; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_370 = 8'h72 == _t_T_2[7:0] ? 8'h40 : _GEN_369; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_371 = 8'h73 == _t_T_2[7:0] ? 8'h8f : _GEN_370; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_372 = 8'h74 == _t_T_2[7:0] ? 8'h92 : _GEN_371; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_373 = 8'h75 == _t_T_2[7:0] ? 8'h9d : _GEN_372; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_374 = 8'h76 == _t_T_2[7:0] ? 8'h38 : _GEN_373; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_375 = 8'h77 == _t_T_2[7:0] ? 8'hf5 : _GEN_374; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_376 = 8'h78 == _t_T_2[7:0] ? 8'hbc : _GEN_375; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_377 = 8'h79 == _t_T_2[7:0] ? 8'hb6 : _GEN_376; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_378 = 8'h7a == _t_T_2[7:0] ? 8'hda : _GEN_377; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_379 = 8'h7b == _t_T_2[7:0] ? 8'h21 : _GEN_378; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_380 = 8'h7c == _t_T_2[7:0] ? 8'h10 : _GEN_379; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_381 = 8'h7d == _t_T_2[7:0] ? 8'hff : _GEN_380; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_382 = 8'h7e == _t_T_2[7:0] ? 8'hf3 : _GEN_381; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_383 = 8'h7f == _t_T_2[7:0] ? 8'hd2 : _GEN_382; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_384 = 8'h80 == _t_T_2[7:0] ? 8'hcd : _GEN_383; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_385 = 8'h81 == _t_T_2[7:0] ? 8'hc : _GEN_384; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_386 = 8'h82 == _t_T_2[7:0] ? 8'h13 : _GEN_385; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_387 = 8'h83 == _t_T_2[7:0] ? 8'hec : _GEN_386; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_388 = 8'h84 == _t_T_2[7:0] ? 8'h5f : _GEN_387; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_389 = 8'h85 == _t_T_2[7:0] ? 8'h97 : _GEN_388; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_390 = 8'h86 == _t_T_2[7:0] ? 8'h44 : _GEN_389; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_391 = 8'h87 == _t_T_2[7:0] ? 8'h17 : _GEN_390; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_392 = 8'h88 == _t_T_2[7:0] ? 8'hc4 : _GEN_391; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_393 = 8'h89 == _t_T_2[7:0] ? 8'ha7 : _GEN_392; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_394 = 8'h8a == _t_T_2[7:0] ? 8'h7e : _GEN_393; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_395 = 8'h8b == _t_T_2[7:0] ? 8'h3d : _GEN_394; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_396 = 8'h8c == _t_T_2[7:0] ? 8'h64 : _GEN_395; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_397 = 8'h8d == _t_T_2[7:0] ? 8'h5d : _GEN_396; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_398 = 8'h8e == _t_T_2[7:0] ? 8'h19 : _GEN_397; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_399 = 8'h8f == _t_T_2[7:0] ? 8'h73 : _GEN_398; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_400 = 8'h90 == _t_T_2[7:0] ? 8'h60 : _GEN_399; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_401 = 8'h91 == _t_T_2[7:0] ? 8'h81 : _GEN_400; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_402 = 8'h92 == _t_T_2[7:0] ? 8'h4f : _GEN_401; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_403 = 8'h93 == _t_T_2[7:0] ? 8'hdc : _GEN_402; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_404 = 8'h94 == _t_T_2[7:0] ? 8'h22 : _GEN_403; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_405 = 8'h95 == _t_T_2[7:0] ? 8'h2a : _GEN_404; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_406 = 8'h96 == _t_T_2[7:0] ? 8'h90 : _GEN_405; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_407 = 8'h97 == _t_T_2[7:0] ? 8'h88 : _GEN_406; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_408 = 8'h98 == _t_T_2[7:0] ? 8'h46 : _GEN_407; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_409 = 8'h99 == _t_T_2[7:0] ? 8'hee : _GEN_408; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_410 = 8'h9a == _t_T_2[7:0] ? 8'hb8 : _GEN_409; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_411 = 8'h9b == _t_T_2[7:0] ? 8'h14 : _GEN_410; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_412 = 8'h9c == _t_T_2[7:0] ? 8'hde : _GEN_411; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_413 = 8'h9d == _t_T_2[7:0] ? 8'h5e : _GEN_412; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_414 = 8'h9e == _t_T_2[7:0] ? 8'hb : _GEN_413; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_415 = 8'h9f == _t_T_2[7:0] ? 8'hdb : _GEN_414; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_416 = 8'ha0 == _t_T_2[7:0] ? 8'he0 : _GEN_415; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_417 = 8'ha1 == _t_T_2[7:0] ? 8'h32 : _GEN_416; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_418 = 8'ha2 == _t_T_2[7:0] ? 8'h3a : _GEN_417; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_419 = 8'ha3 == _t_T_2[7:0] ? 8'ha : _GEN_418; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_420 = 8'ha4 == _t_T_2[7:0] ? 8'h49 : _GEN_419; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_421 = 8'ha5 == _t_T_2[7:0] ? 8'h6 : _GEN_420; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_422 = 8'ha6 == _t_T_2[7:0] ? 8'h24 : _GEN_421; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_423 = 8'ha7 == _t_T_2[7:0] ? 8'h5c : _GEN_422; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_424 = 8'ha8 == _t_T_2[7:0] ? 8'hc2 : _GEN_423; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_425 = 8'ha9 == _t_T_2[7:0] ? 8'hd3 : _GEN_424; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_426 = 8'haa == _t_T_2[7:0] ? 8'hac : _GEN_425; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_427 = 8'hab == _t_T_2[7:0] ? 8'h62 : _GEN_426; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_428 = 8'hac == _t_T_2[7:0] ? 8'h91 : _GEN_427; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_429 = 8'had == _t_T_2[7:0] ? 8'h95 : _GEN_428; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_430 = 8'hae == _t_T_2[7:0] ? 8'he4 : _GEN_429; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_431 = 8'haf == _t_T_2[7:0] ? 8'h79 : _GEN_430; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_432 = 8'hb0 == _t_T_2[7:0] ? 8'he7 : _GEN_431; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_433 = 8'hb1 == _t_T_2[7:0] ? 8'hc8 : _GEN_432; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_434 = 8'hb2 == _t_T_2[7:0] ? 8'h37 : _GEN_433; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_435 = 8'hb3 == _t_T_2[7:0] ? 8'h6d : _GEN_434; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_436 = 8'hb4 == _t_T_2[7:0] ? 8'h8d : _GEN_435; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_437 = 8'hb5 == _t_T_2[7:0] ? 8'hd5 : _GEN_436; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_438 = 8'hb6 == _t_T_2[7:0] ? 8'h4e : _GEN_437; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_439 = 8'hb7 == _t_T_2[7:0] ? 8'ha9 : _GEN_438; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_440 = 8'hb8 == _t_T_2[7:0] ? 8'h6c : _GEN_439; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_441 = 8'hb9 == _t_T_2[7:0] ? 8'h56 : _GEN_440; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_442 = 8'hba == _t_T_2[7:0] ? 8'hf4 : _GEN_441; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_443 = 8'hbb == _t_T_2[7:0] ? 8'hea : _GEN_442; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_444 = 8'hbc == _t_T_2[7:0] ? 8'h65 : _GEN_443; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_445 = 8'hbd == _t_T_2[7:0] ? 8'h7a : _GEN_444; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_446 = 8'hbe == _t_T_2[7:0] ? 8'hae : _GEN_445; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_447 = 8'hbf == _t_T_2[7:0] ? 8'h8 : _GEN_446; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_448 = 8'hc0 == _t_T_2[7:0] ? 8'hba : _GEN_447; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_449 = 8'hc1 == _t_T_2[7:0] ? 8'h78 : _GEN_448; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_450 = 8'hc2 == _t_T_2[7:0] ? 8'h25 : _GEN_449; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_451 = 8'hc3 == _t_T_2[7:0] ? 8'h2e : _GEN_450; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_452 = 8'hc4 == _t_T_2[7:0] ? 8'h1c : _GEN_451; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_453 = 8'hc5 == _t_T_2[7:0] ? 8'ha6 : _GEN_452; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_454 = 8'hc6 == _t_T_2[7:0] ? 8'hb4 : _GEN_453; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_455 = 8'hc7 == _t_T_2[7:0] ? 8'hc6 : _GEN_454; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_456 = 8'hc8 == _t_T_2[7:0] ? 8'he8 : _GEN_455; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_457 = 8'hc9 == _t_T_2[7:0] ? 8'hdd : _GEN_456; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_458 = 8'hca == _t_T_2[7:0] ? 8'h74 : _GEN_457; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_459 = 8'hcb == _t_T_2[7:0] ? 8'h1f : _GEN_458; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_460 = 8'hcc == _t_T_2[7:0] ? 8'h4b : _GEN_459; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_461 = 8'hcd == _t_T_2[7:0] ? 8'hbd : _GEN_460; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_462 = 8'hce == _t_T_2[7:0] ? 8'h8b : _GEN_461; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_463 = 8'hcf == _t_T_2[7:0] ? 8'h8a : _GEN_462; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_464 = 8'hd0 == _t_T_2[7:0] ? 8'h70 : _GEN_463; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_465 = 8'hd1 == _t_T_2[7:0] ? 8'h3e : _GEN_464; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_466 = 8'hd2 == _t_T_2[7:0] ? 8'hb5 : _GEN_465; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_467 = 8'hd3 == _t_T_2[7:0] ? 8'h66 : _GEN_466; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_468 = 8'hd4 == _t_T_2[7:0] ? 8'h48 : _GEN_467; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_469 = 8'hd5 == _t_T_2[7:0] ? 8'h3 : _GEN_468; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_470 = 8'hd6 == _t_T_2[7:0] ? 8'hf6 : _GEN_469; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_471 = 8'hd7 == _t_T_2[7:0] ? 8'he : _GEN_470; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_472 = 8'hd8 == _t_T_2[7:0] ? 8'h61 : _GEN_471; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_473 = 8'hd9 == _t_T_2[7:0] ? 8'h35 : _GEN_472; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_474 = 8'hda == _t_T_2[7:0] ? 8'h57 : _GEN_473; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_475 = 8'hdb == _t_T_2[7:0] ? 8'hb9 : _GEN_474; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_476 = 8'hdc == _t_T_2[7:0] ? 8'h86 : _GEN_475; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_477 = 8'hdd == _t_T_2[7:0] ? 8'hc1 : _GEN_476; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_478 = 8'hde == _t_T_2[7:0] ? 8'h1d : _GEN_477; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_479 = 8'hdf == _t_T_2[7:0] ? 8'h9e : _GEN_478; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_480 = 8'he0 == _t_T_2[7:0] ? 8'he1 : _GEN_479; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_481 = 8'he1 == _t_T_2[7:0] ? 8'hf8 : _GEN_480; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_482 = 8'he2 == _t_T_2[7:0] ? 8'h98 : _GEN_481; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_483 = 8'he3 == _t_T_2[7:0] ? 8'h11 : _GEN_482; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_484 = 8'he4 == _t_T_2[7:0] ? 8'h69 : _GEN_483; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_485 = 8'he5 == _t_T_2[7:0] ? 8'hd9 : _GEN_484; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_486 = 8'he6 == _t_T_2[7:0] ? 8'h8e : _GEN_485; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_487 = 8'he7 == _t_T_2[7:0] ? 8'h94 : _GEN_486; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_488 = 8'he8 == _t_T_2[7:0] ? 8'h9b : _GEN_487; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_489 = 8'he9 == _t_T_2[7:0] ? 8'h1e : _GEN_488; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_490 = 8'hea == _t_T_2[7:0] ? 8'h87 : _GEN_489; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_491 = 8'heb == _t_T_2[7:0] ? 8'he9 : _GEN_490; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_492 = 8'hec == _t_T_2[7:0] ? 8'hce : _GEN_491; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_493 = 8'hed == _t_T_2[7:0] ? 8'h55 : _GEN_492; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_494 = 8'hee == _t_T_2[7:0] ? 8'h28 : _GEN_493; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_495 = 8'hef == _t_T_2[7:0] ? 8'hdf : _GEN_494; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_496 = 8'hf0 == _t_T_2[7:0] ? 8'h8c : _GEN_495; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_497 = 8'hf1 == _t_T_2[7:0] ? 8'ha1 : _GEN_496; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_498 = 8'hf2 == _t_T_2[7:0] ? 8'h89 : _GEN_497; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_499 = 8'hf3 == _t_T_2[7:0] ? 8'hd : _GEN_498; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_500 = 8'hf4 == _t_T_2[7:0] ? 8'hbf : _GEN_499; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_501 = 8'hf5 == _t_T_2[7:0] ? 8'he6 : _GEN_500; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_502 = 8'hf6 == _t_T_2[7:0] ? 8'h42 : _GEN_501; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_503 = 8'hf7 == _t_T_2[7:0] ? 8'h68 : _GEN_502; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_504 = 8'hf8 == _t_T_2[7:0] ? 8'h41 : _GEN_503; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_505 = 8'hf9 == _t_T_2[7:0] ? 8'h99 : _GEN_504; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_506 = 8'hfa == _t_T_2[7:0] ? 8'h2d : _GEN_505; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_507 = 8'hfb == _t_T_2[7:0] ? 8'hf : _GEN_506; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_508 = 8'hfc == _t_T_2[7:0] ? 8'hb0 : _GEN_507; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_509 = 8'hfd == _t_T_2[7:0] ? 8'h54 : _GEN_508; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_510 = 8'hfe == _t_T_2[7:0] ? 8'hbb : _GEN_509; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_511 = 8'hff == _t_T_2[7:0] ? 8'h16 : _GEN_510; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_513 = 8'h1 == _t_T_2[31:24] ? 8'h7c : 8'h63; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_514 = 8'h2 == _t_T_2[31:24] ? 8'h77 : _GEN_513; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_515 = 8'h3 == _t_T_2[31:24] ? 8'h7b : _GEN_514; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_516 = 8'h4 == _t_T_2[31:24] ? 8'hf2 : _GEN_515; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_517 = 8'h5 == _t_T_2[31:24] ? 8'h6b : _GEN_516; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_518 = 8'h6 == _t_T_2[31:24] ? 8'h6f : _GEN_517; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_519 = 8'h7 == _t_T_2[31:24] ? 8'hc5 : _GEN_518; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_520 = 8'h8 == _t_T_2[31:24] ? 8'h30 : _GEN_519; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_521 = 8'h9 == _t_T_2[31:24] ? 8'h1 : _GEN_520; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_522 = 8'ha == _t_T_2[31:24] ? 8'h67 : _GEN_521; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_523 = 8'hb == _t_T_2[31:24] ? 8'h2b : _GEN_522; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_524 = 8'hc == _t_T_2[31:24] ? 8'hfe : _GEN_523; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_525 = 8'hd == _t_T_2[31:24] ? 8'hd7 : _GEN_524; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_526 = 8'he == _t_T_2[31:24] ? 8'hab : _GEN_525; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_527 = 8'hf == _t_T_2[31:24] ? 8'h76 : _GEN_526; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_528 = 8'h10 == _t_T_2[31:24] ? 8'hca : _GEN_527; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_529 = 8'h11 == _t_T_2[31:24] ? 8'h82 : _GEN_528; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_530 = 8'h12 == _t_T_2[31:24] ? 8'hc9 : _GEN_529; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_531 = 8'h13 == _t_T_2[31:24] ? 8'h7d : _GEN_530; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_532 = 8'h14 == _t_T_2[31:24] ? 8'hfa : _GEN_531; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_533 = 8'h15 == _t_T_2[31:24] ? 8'h59 : _GEN_532; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_534 = 8'h16 == _t_T_2[31:24] ? 8'h47 : _GEN_533; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_535 = 8'h17 == _t_T_2[31:24] ? 8'hf0 : _GEN_534; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_536 = 8'h18 == _t_T_2[31:24] ? 8'had : _GEN_535; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_537 = 8'h19 == _t_T_2[31:24] ? 8'hd4 : _GEN_536; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_538 = 8'h1a == _t_T_2[31:24] ? 8'ha2 : _GEN_537; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_539 = 8'h1b == _t_T_2[31:24] ? 8'haf : _GEN_538; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_540 = 8'h1c == _t_T_2[31:24] ? 8'h9c : _GEN_539; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_541 = 8'h1d == _t_T_2[31:24] ? 8'ha4 : _GEN_540; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_542 = 8'h1e == _t_T_2[31:24] ? 8'h72 : _GEN_541; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_543 = 8'h1f == _t_T_2[31:24] ? 8'hc0 : _GEN_542; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_544 = 8'h20 == _t_T_2[31:24] ? 8'hb7 : _GEN_543; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_545 = 8'h21 == _t_T_2[31:24] ? 8'hfd : _GEN_544; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_546 = 8'h22 == _t_T_2[31:24] ? 8'h93 : _GEN_545; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_547 = 8'h23 == _t_T_2[31:24] ? 8'h26 : _GEN_546; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_548 = 8'h24 == _t_T_2[31:24] ? 8'h36 : _GEN_547; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_549 = 8'h25 == _t_T_2[31:24] ? 8'h3f : _GEN_548; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_550 = 8'h26 == _t_T_2[31:24] ? 8'hf7 : _GEN_549; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_551 = 8'h27 == _t_T_2[31:24] ? 8'hcc : _GEN_550; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_552 = 8'h28 == _t_T_2[31:24] ? 8'h34 : _GEN_551; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_553 = 8'h29 == _t_T_2[31:24] ? 8'ha5 : _GEN_552; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_554 = 8'h2a == _t_T_2[31:24] ? 8'he5 : _GEN_553; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_555 = 8'h2b == _t_T_2[31:24] ? 8'hf1 : _GEN_554; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_556 = 8'h2c == _t_T_2[31:24] ? 8'h71 : _GEN_555; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_557 = 8'h2d == _t_T_2[31:24] ? 8'hd8 : _GEN_556; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_558 = 8'h2e == _t_T_2[31:24] ? 8'h31 : _GEN_557; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_559 = 8'h2f == _t_T_2[31:24] ? 8'h15 : _GEN_558; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_560 = 8'h30 == _t_T_2[31:24] ? 8'h4 : _GEN_559; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_561 = 8'h31 == _t_T_2[31:24] ? 8'hc7 : _GEN_560; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_562 = 8'h32 == _t_T_2[31:24] ? 8'h23 : _GEN_561; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_563 = 8'h33 == _t_T_2[31:24] ? 8'hc3 : _GEN_562; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_564 = 8'h34 == _t_T_2[31:24] ? 8'h18 : _GEN_563; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_565 = 8'h35 == _t_T_2[31:24] ? 8'h96 : _GEN_564; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_566 = 8'h36 == _t_T_2[31:24] ? 8'h5 : _GEN_565; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_567 = 8'h37 == _t_T_2[31:24] ? 8'h9a : _GEN_566; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_568 = 8'h38 == _t_T_2[31:24] ? 8'h7 : _GEN_567; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_569 = 8'h39 == _t_T_2[31:24] ? 8'h12 : _GEN_568; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_570 = 8'h3a == _t_T_2[31:24] ? 8'h80 : _GEN_569; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_571 = 8'h3b == _t_T_2[31:24] ? 8'he2 : _GEN_570; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_572 = 8'h3c == _t_T_2[31:24] ? 8'heb : _GEN_571; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_573 = 8'h3d == _t_T_2[31:24] ? 8'h27 : _GEN_572; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_574 = 8'h3e == _t_T_2[31:24] ? 8'hb2 : _GEN_573; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_575 = 8'h3f == _t_T_2[31:24] ? 8'h75 : _GEN_574; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_576 = 8'h40 == _t_T_2[31:24] ? 8'h9 : _GEN_575; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_577 = 8'h41 == _t_T_2[31:24] ? 8'h83 : _GEN_576; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_578 = 8'h42 == _t_T_2[31:24] ? 8'h2c : _GEN_577; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_579 = 8'h43 == _t_T_2[31:24] ? 8'h1a : _GEN_578; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_580 = 8'h44 == _t_T_2[31:24] ? 8'h1b : _GEN_579; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_581 = 8'h45 == _t_T_2[31:24] ? 8'h6e : _GEN_580; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_582 = 8'h46 == _t_T_2[31:24] ? 8'h5a : _GEN_581; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_583 = 8'h47 == _t_T_2[31:24] ? 8'ha0 : _GEN_582; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_584 = 8'h48 == _t_T_2[31:24] ? 8'h52 : _GEN_583; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_585 = 8'h49 == _t_T_2[31:24] ? 8'h3b : _GEN_584; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_586 = 8'h4a == _t_T_2[31:24] ? 8'hd6 : _GEN_585; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_587 = 8'h4b == _t_T_2[31:24] ? 8'hb3 : _GEN_586; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_588 = 8'h4c == _t_T_2[31:24] ? 8'h29 : _GEN_587; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_589 = 8'h4d == _t_T_2[31:24] ? 8'he3 : _GEN_588; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_590 = 8'h4e == _t_T_2[31:24] ? 8'h2f : _GEN_589; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_591 = 8'h4f == _t_T_2[31:24] ? 8'h84 : _GEN_590; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_592 = 8'h50 == _t_T_2[31:24] ? 8'h53 : _GEN_591; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_593 = 8'h51 == _t_T_2[31:24] ? 8'hd1 : _GEN_592; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_594 = 8'h52 == _t_T_2[31:24] ? 8'h0 : _GEN_593; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_595 = 8'h53 == _t_T_2[31:24] ? 8'hed : _GEN_594; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_596 = 8'h54 == _t_T_2[31:24] ? 8'h20 : _GEN_595; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_597 = 8'h55 == _t_T_2[31:24] ? 8'hfc : _GEN_596; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_598 = 8'h56 == _t_T_2[31:24] ? 8'hb1 : _GEN_597; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_599 = 8'h57 == _t_T_2[31:24] ? 8'h5b : _GEN_598; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_600 = 8'h58 == _t_T_2[31:24] ? 8'h6a : _GEN_599; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_601 = 8'h59 == _t_T_2[31:24] ? 8'hcb : _GEN_600; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_602 = 8'h5a == _t_T_2[31:24] ? 8'hbe : _GEN_601; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_603 = 8'h5b == _t_T_2[31:24] ? 8'h39 : _GEN_602; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_604 = 8'h5c == _t_T_2[31:24] ? 8'h4a : _GEN_603; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_605 = 8'h5d == _t_T_2[31:24] ? 8'h4c : _GEN_604; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_606 = 8'h5e == _t_T_2[31:24] ? 8'h58 : _GEN_605; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_607 = 8'h5f == _t_T_2[31:24] ? 8'hcf : _GEN_606; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_608 = 8'h60 == _t_T_2[31:24] ? 8'hd0 : _GEN_607; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_609 = 8'h61 == _t_T_2[31:24] ? 8'hef : _GEN_608; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_610 = 8'h62 == _t_T_2[31:24] ? 8'haa : _GEN_609; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_611 = 8'h63 == _t_T_2[31:24] ? 8'hfb : _GEN_610; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_612 = 8'h64 == _t_T_2[31:24] ? 8'h43 : _GEN_611; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_613 = 8'h65 == _t_T_2[31:24] ? 8'h4d : _GEN_612; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_614 = 8'h66 == _t_T_2[31:24] ? 8'h33 : _GEN_613; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_615 = 8'h67 == _t_T_2[31:24] ? 8'h85 : _GEN_614; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_616 = 8'h68 == _t_T_2[31:24] ? 8'h45 : _GEN_615; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_617 = 8'h69 == _t_T_2[31:24] ? 8'hf9 : _GEN_616; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_618 = 8'h6a == _t_T_2[31:24] ? 8'h2 : _GEN_617; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_619 = 8'h6b == _t_T_2[31:24] ? 8'h7f : _GEN_618; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_620 = 8'h6c == _t_T_2[31:24] ? 8'h50 : _GEN_619; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_621 = 8'h6d == _t_T_2[31:24] ? 8'h3c : _GEN_620; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_622 = 8'h6e == _t_T_2[31:24] ? 8'h9f : _GEN_621; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_623 = 8'h6f == _t_T_2[31:24] ? 8'ha8 : _GEN_622; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_624 = 8'h70 == _t_T_2[31:24] ? 8'h51 : _GEN_623; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_625 = 8'h71 == _t_T_2[31:24] ? 8'ha3 : _GEN_624; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_626 = 8'h72 == _t_T_2[31:24] ? 8'h40 : _GEN_625; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_627 = 8'h73 == _t_T_2[31:24] ? 8'h8f : _GEN_626; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_628 = 8'h74 == _t_T_2[31:24] ? 8'h92 : _GEN_627; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_629 = 8'h75 == _t_T_2[31:24] ? 8'h9d : _GEN_628; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_630 = 8'h76 == _t_T_2[31:24] ? 8'h38 : _GEN_629; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_631 = 8'h77 == _t_T_2[31:24] ? 8'hf5 : _GEN_630; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_632 = 8'h78 == _t_T_2[31:24] ? 8'hbc : _GEN_631; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_633 = 8'h79 == _t_T_2[31:24] ? 8'hb6 : _GEN_632; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_634 = 8'h7a == _t_T_2[31:24] ? 8'hda : _GEN_633; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_635 = 8'h7b == _t_T_2[31:24] ? 8'h21 : _GEN_634; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_636 = 8'h7c == _t_T_2[31:24] ? 8'h10 : _GEN_635; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_637 = 8'h7d == _t_T_2[31:24] ? 8'hff : _GEN_636; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_638 = 8'h7e == _t_T_2[31:24] ? 8'hf3 : _GEN_637; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_639 = 8'h7f == _t_T_2[31:24] ? 8'hd2 : _GEN_638; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_640 = 8'h80 == _t_T_2[31:24] ? 8'hcd : _GEN_639; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_641 = 8'h81 == _t_T_2[31:24] ? 8'hc : _GEN_640; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_642 = 8'h82 == _t_T_2[31:24] ? 8'h13 : _GEN_641; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_643 = 8'h83 == _t_T_2[31:24] ? 8'hec : _GEN_642; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_644 = 8'h84 == _t_T_2[31:24] ? 8'h5f : _GEN_643; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_645 = 8'h85 == _t_T_2[31:24] ? 8'h97 : _GEN_644; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_646 = 8'h86 == _t_T_2[31:24] ? 8'h44 : _GEN_645; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_647 = 8'h87 == _t_T_2[31:24] ? 8'h17 : _GEN_646; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_648 = 8'h88 == _t_T_2[31:24] ? 8'hc4 : _GEN_647; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_649 = 8'h89 == _t_T_2[31:24] ? 8'ha7 : _GEN_648; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_650 = 8'h8a == _t_T_2[31:24] ? 8'h7e : _GEN_649; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_651 = 8'h8b == _t_T_2[31:24] ? 8'h3d : _GEN_650; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_652 = 8'h8c == _t_T_2[31:24] ? 8'h64 : _GEN_651; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_653 = 8'h8d == _t_T_2[31:24] ? 8'h5d : _GEN_652; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_654 = 8'h8e == _t_T_2[31:24] ? 8'h19 : _GEN_653; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_655 = 8'h8f == _t_T_2[31:24] ? 8'h73 : _GEN_654; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_656 = 8'h90 == _t_T_2[31:24] ? 8'h60 : _GEN_655; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_657 = 8'h91 == _t_T_2[31:24] ? 8'h81 : _GEN_656; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_658 = 8'h92 == _t_T_2[31:24] ? 8'h4f : _GEN_657; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_659 = 8'h93 == _t_T_2[31:24] ? 8'hdc : _GEN_658; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_660 = 8'h94 == _t_T_2[31:24] ? 8'h22 : _GEN_659; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_661 = 8'h95 == _t_T_2[31:24] ? 8'h2a : _GEN_660; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_662 = 8'h96 == _t_T_2[31:24] ? 8'h90 : _GEN_661; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_663 = 8'h97 == _t_T_2[31:24] ? 8'h88 : _GEN_662; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_664 = 8'h98 == _t_T_2[31:24] ? 8'h46 : _GEN_663; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_665 = 8'h99 == _t_T_2[31:24] ? 8'hee : _GEN_664; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_666 = 8'h9a == _t_T_2[31:24] ? 8'hb8 : _GEN_665; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_667 = 8'h9b == _t_T_2[31:24] ? 8'h14 : _GEN_666; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_668 = 8'h9c == _t_T_2[31:24] ? 8'hde : _GEN_667; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_669 = 8'h9d == _t_T_2[31:24] ? 8'h5e : _GEN_668; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_670 = 8'h9e == _t_T_2[31:24] ? 8'hb : _GEN_669; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_671 = 8'h9f == _t_T_2[31:24] ? 8'hdb : _GEN_670; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_672 = 8'ha0 == _t_T_2[31:24] ? 8'he0 : _GEN_671; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_673 = 8'ha1 == _t_T_2[31:24] ? 8'h32 : _GEN_672; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_674 = 8'ha2 == _t_T_2[31:24] ? 8'h3a : _GEN_673; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_675 = 8'ha3 == _t_T_2[31:24] ? 8'ha : _GEN_674; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_676 = 8'ha4 == _t_T_2[31:24] ? 8'h49 : _GEN_675; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_677 = 8'ha5 == _t_T_2[31:24] ? 8'h6 : _GEN_676; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_678 = 8'ha6 == _t_T_2[31:24] ? 8'h24 : _GEN_677; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_679 = 8'ha7 == _t_T_2[31:24] ? 8'h5c : _GEN_678; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_680 = 8'ha8 == _t_T_2[31:24] ? 8'hc2 : _GEN_679; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_681 = 8'ha9 == _t_T_2[31:24] ? 8'hd3 : _GEN_680; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_682 = 8'haa == _t_T_2[31:24] ? 8'hac : _GEN_681; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_683 = 8'hab == _t_T_2[31:24] ? 8'h62 : _GEN_682; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_684 = 8'hac == _t_T_2[31:24] ? 8'h91 : _GEN_683; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_685 = 8'had == _t_T_2[31:24] ? 8'h95 : _GEN_684; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_686 = 8'hae == _t_T_2[31:24] ? 8'he4 : _GEN_685; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_687 = 8'haf == _t_T_2[31:24] ? 8'h79 : _GEN_686; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_688 = 8'hb0 == _t_T_2[31:24] ? 8'he7 : _GEN_687; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_689 = 8'hb1 == _t_T_2[31:24] ? 8'hc8 : _GEN_688; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_690 = 8'hb2 == _t_T_2[31:24] ? 8'h37 : _GEN_689; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_691 = 8'hb3 == _t_T_2[31:24] ? 8'h6d : _GEN_690; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_692 = 8'hb4 == _t_T_2[31:24] ? 8'h8d : _GEN_691; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_693 = 8'hb5 == _t_T_2[31:24] ? 8'hd5 : _GEN_692; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_694 = 8'hb6 == _t_T_2[31:24] ? 8'h4e : _GEN_693; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_695 = 8'hb7 == _t_T_2[31:24] ? 8'ha9 : _GEN_694; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_696 = 8'hb8 == _t_T_2[31:24] ? 8'h6c : _GEN_695; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_697 = 8'hb9 == _t_T_2[31:24] ? 8'h56 : _GEN_696; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_698 = 8'hba == _t_T_2[31:24] ? 8'hf4 : _GEN_697; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_699 = 8'hbb == _t_T_2[31:24] ? 8'hea : _GEN_698; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_700 = 8'hbc == _t_T_2[31:24] ? 8'h65 : _GEN_699; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_701 = 8'hbd == _t_T_2[31:24] ? 8'h7a : _GEN_700; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_702 = 8'hbe == _t_T_2[31:24] ? 8'hae : _GEN_701; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_703 = 8'hbf == _t_T_2[31:24] ? 8'h8 : _GEN_702; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_704 = 8'hc0 == _t_T_2[31:24] ? 8'hba : _GEN_703; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_705 = 8'hc1 == _t_T_2[31:24] ? 8'h78 : _GEN_704; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_706 = 8'hc2 == _t_T_2[31:24] ? 8'h25 : _GEN_705; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_707 = 8'hc3 == _t_T_2[31:24] ? 8'h2e : _GEN_706; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_708 = 8'hc4 == _t_T_2[31:24] ? 8'h1c : _GEN_707; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_709 = 8'hc5 == _t_T_2[31:24] ? 8'ha6 : _GEN_708; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_710 = 8'hc6 == _t_T_2[31:24] ? 8'hb4 : _GEN_709; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_711 = 8'hc7 == _t_T_2[31:24] ? 8'hc6 : _GEN_710; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_712 = 8'hc8 == _t_T_2[31:24] ? 8'he8 : _GEN_711; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_713 = 8'hc9 == _t_T_2[31:24] ? 8'hdd : _GEN_712; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_714 = 8'hca == _t_T_2[31:24] ? 8'h74 : _GEN_713; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_715 = 8'hcb == _t_T_2[31:24] ? 8'h1f : _GEN_714; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_716 = 8'hcc == _t_T_2[31:24] ? 8'h4b : _GEN_715; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_717 = 8'hcd == _t_T_2[31:24] ? 8'hbd : _GEN_716; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_718 = 8'hce == _t_T_2[31:24] ? 8'h8b : _GEN_717; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_719 = 8'hcf == _t_T_2[31:24] ? 8'h8a : _GEN_718; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_720 = 8'hd0 == _t_T_2[31:24] ? 8'h70 : _GEN_719; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_721 = 8'hd1 == _t_T_2[31:24] ? 8'h3e : _GEN_720; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_722 = 8'hd2 == _t_T_2[31:24] ? 8'hb5 : _GEN_721; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_723 = 8'hd3 == _t_T_2[31:24] ? 8'h66 : _GEN_722; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_724 = 8'hd4 == _t_T_2[31:24] ? 8'h48 : _GEN_723; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_725 = 8'hd5 == _t_T_2[31:24] ? 8'h3 : _GEN_724; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_726 = 8'hd6 == _t_T_2[31:24] ? 8'hf6 : _GEN_725; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_727 = 8'hd7 == _t_T_2[31:24] ? 8'he : _GEN_726; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_728 = 8'hd8 == _t_T_2[31:24] ? 8'h61 : _GEN_727; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_729 = 8'hd9 == _t_T_2[31:24] ? 8'h35 : _GEN_728; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_730 = 8'hda == _t_T_2[31:24] ? 8'h57 : _GEN_729; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_731 = 8'hdb == _t_T_2[31:24] ? 8'hb9 : _GEN_730; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_732 = 8'hdc == _t_T_2[31:24] ? 8'h86 : _GEN_731; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_733 = 8'hdd == _t_T_2[31:24] ? 8'hc1 : _GEN_732; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_734 = 8'hde == _t_T_2[31:24] ? 8'h1d : _GEN_733; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_735 = 8'hdf == _t_T_2[31:24] ? 8'h9e : _GEN_734; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_736 = 8'he0 == _t_T_2[31:24] ? 8'he1 : _GEN_735; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_737 = 8'he1 == _t_T_2[31:24] ? 8'hf8 : _GEN_736; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_738 = 8'he2 == _t_T_2[31:24] ? 8'h98 : _GEN_737; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_739 = 8'he3 == _t_T_2[31:24] ? 8'h11 : _GEN_738; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_740 = 8'he4 == _t_T_2[31:24] ? 8'h69 : _GEN_739; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_741 = 8'he5 == _t_T_2[31:24] ? 8'hd9 : _GEN_740; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_742 = 8'he6 == _t_T_2[31:24] ? 8'h8e : _GEN_741; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_743 = 8'he7 == _t_T_2[31:24] ? 8'h94 : _GEN_742; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_744 = 8'he8 == _t_T_2[31:24] ? 8'h9b : _GEN_743; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_745 = 8'he9 == _t_T_2[31:24] ? 8'h1e : _GEN_744; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_746 = 8'hea == _t_T_2[31:24] ? 8'h87 : _GEN_745; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_747 = 8'heb == _t_T_2[31:24] ? 8'he9 : _GEN_746; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_748 = 8'hec == _t_T_2[31:24] ? 8'hce : _GEN_747; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_749 = 8'hed == _t_T_2[31:24] ? 8'h55 : _GEN_748; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_750 = 8'hee == _t_T_2[31:24] ? 8'h28 : _GEN_749; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_751 = 8'hef == _t_T_2[31:24] ? 8'hdf : _GEN_750; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_752 = 8'hf0 == _t_T_2[31:24] ? 8'h8c : _GEN_751; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_753 = 8'hf1 == _t_T_2[31:24] ? 8'ha1 : _GEN_752; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_754 = 8'hf2 == _t_T_2[31:24] ? 8'h89 : _GEN_753; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_755 = 8'hf3 == _t_T_2[31:24] ? 8'hd : _GEN_754; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_756 = 8'hf4 == _t_T_2[31:24] ? 8'hbf : _GEN_755; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_757 = 8'hf5 == _t_T_2[31:24] ? 8'he6 : _GEN_756; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_758 = 8'hf6 == _t_T_2[31:24] ? 8'h42 : _GEN_757; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_759 = 8'hf7 == _t_T_2[31:24] ? 8'h68 : _GEN_758; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_760 = 8'hf8 == _t_T_2[31:24] ? 8'h41 : _GEN_759; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_761 = 8'hf9 == _t_T_2[31:24] ? 8'h99 : _GEN_760; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_762 = 8'hfa == _t_T_2[31:24] ? 8'h2d : _GEN_761; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_763 = 8'hfb == _t_T_2[31:24] ? 8'hf : _GEN_762; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_764 = 8'hfc == _t_T_2[31:24] ? 8'hb0 : _GEN_763; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_765 = 8'hfd == _t_T_2[31:24] ? 8'h54 : _GEN_764; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_766 = 8'hfe == _t_T_2[31:24] ? 8'hbb : _GEN_765; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_767 = 8'hff == _t_T_2[31:24] ? 8'h16 : _GEN_766; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_769 = 8'h1 == _t_T_2[23:16] ? 8'h7c : 8'h63; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_770 = 8'h2 == _t_T_2[23:16] ? 8'h77 : _GEN_769; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_771 = 8'h3 == _t_T_2[23:16] ? 8'h7b : _GEN_770; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_772 = 8'h4 == _t_T_2[23:16] ? 8'hf2 : _GEN_771; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_773 = 8'h5 == _t_T_2[23:16] ? 8'h6b : _GEN_772; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_774 = 8'h6 == _t_T_2[23:16] ? 8'h6f : _GEN_773; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_775 = 8'h7 == _t_T_2[23:16] ? 8'hc5 : _GEN_774; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_776 = 8'h8 == _t_T_2[23:16] ? 8'h30 : _GEN_775; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_777 = 8'h9 == _t_T_2[23:16] ? 8'h1 : _GEN_776; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_778 = 8'ha == _t_T_2[23:16] ? 8'h67 : _GEN_777; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_779 = 8'hb == _t_T_2[23:16] ? 8'h2b : _GEN_778; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_780 = 8'hc == _t_T_2[23:16] ? 8'hfe : _GEN_779; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_781 = 8'hd == _t_T_2[23:16] ? 8'hd7 : _GEN_780; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_782 = 8'he == _t_T_2[23:16] ? 8'hab : _GEN_781; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_783 = 8'hf == _t_T_2[23:16] ? 8'h76 : _GEN_782; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_784 = 8'h10 == _t_T_2[23:16] ? 8'hca : _GEN_783; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_785 = 8'h11 == _t_T_2[23:16] ? 8'h82 : _GEN_784; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_786 = 8'h12 == _t_T_2[23:16] ? 8'hc9 : _GEN_785; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_787 = 8'h13 == _t_T_2[23:16] ? 8'h7d : _GEN_786; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_788 = 8'h14 == _t_T_2[23:16] ? 8'hfa : _GEN_787; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_789 = 8'h15 == _t_T_2[23:16] ? 8'h59 : _GEN_788; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_790 = 8'h16 == _t_T_2[23:16] ? 8'h47 : _GEN_789; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_791 = 8'h17 == _t_T_2[23:16] ? 8'hf0 : _GEN_790; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_792 = 8'h18 == _t_T_2[23:16] ? 8'had : _GEN_791; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_793 = 8'h19 == _t_T_2[23:16] ? 8'hd4 : _GEN_792; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_794 = 8'h1a == _t_T_2[23:16] ? 8'ha2 : _GEN_793; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_795 = 8'h1b == _t_T_2[23:16] ? 8'haf : _GEN_794; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_796 = 8'h1c == _t_T_2[23:16] ? 8'h9c : _GEN_795; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_797 = 8'h1d == _t_T_2[23:16] ? 8'ha4 : _GEN_796; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_798 = 8'h1e == _t_T_2[23:16] ? 8'h72 : _GEN_797; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_799 = 8'h1f == _t_T_2[23:16] ? 8'hc0 : _GEN_798; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_800 = 8'h20 == _t_T_2[23:16] ? 8'hb7 : _GEN_799; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_801 = 8'h21 == _t_T_2[23:16] ? 8'hfd : _GEN_800; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_802 = 8'h22 == _t_T_2[23:16] ? 8'h93 : _GEN_801; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_803 = 8'h23 == _t_T_2[23:16] ? 8'h26 : _GEN_802; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_804 = 8'h24 == _t_T_2[23:16] ? 8'h36 : _GEN_803; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_805 = 8'h25 == _t_T_2[23:16] ? 8'h3f : _GEN_804; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_806 = 8'h26 == _t_T_2[23:16] ? 8'hf7 : _GEN_805; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_807 = 8'h27 == _t_T_2[23:16] ? 8'hcc : _GEN_806; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_808 = 8'h28 == _t_T_2[23:16] ? 8'h34 : _GEN_807; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_809 = 8'h29 == _t_T_2[23:16] ? 8'ha5 : _GEN_808; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_810 = 8'h2a == _t_T_2[23:16] ? 8'he5 : _GEN_809; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_811 = 8'h2b == _t_T_2[23:16] ? 8'hf1 : _GEN_810; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_812 = 8'h2c == _t_T_2[23:16] ? 8'h71 : _GEN_811; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_813 = 8'h2d == _t_T_2[23:16] ? 8'hd8 : _GEN_812; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_814 = 8'h2e == _t_T_2[23:16] ? 8'h31 : _GEN_813; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_815 = 8'h2f == _t_T_2[23:16] ? 8'h15 : _GEN_814; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_816 = 8'h30 == _t_T_2[23:16] ? 8'h4 : _GEN_815; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_817 = 8'h31 == _t_T_2[23:16] ? 8'hc7 : _GEN_816; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_818 = 8'h32 == _t_T_2[23:16] ? 8'h23 : _GEN_817; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_819 = 8'h33 == _t_T_2[23:16] ? 8'hc3 : _GEN_818; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_820 = 8'h34 == _t_T_2[23:16] ? 8'h18 : _GEN_819; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_821 = 8'h35 == _t_T_2[23:16] ? 8'h96 : _GEN_820; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_822 = 8'h36 == _t_T_2[23:16] ? 8'h5 : _GEN_821; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_823 = 8'h37 == _t_T_2[23:16] ? 8'h9a : _GEN_822; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_824 = 8'h38 == _t_T_2[23:16] ? 8'h7 : _GEN_823; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_825 = 8'h39 == _t_T_2[23:16] ? 8'h12 : _GEN_824; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_826 = 8'h3a == _t_T_2[23:16] ? 8'h80 : _GEN_825; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_827 = 8'h3b == _t_T_2[23:16] ? 8'he2 : _GEN_826; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_828 = 8'h3c == _t_T_2[23:16] ? 8'heb : _GEN_827; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_829 = 8'h3d == _t_T_2[23:16] ? 8'h27 : _GEN_828; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_830 = 8'h3e == _t_T_2[23:16] ? 8'hb2 : _GEN_829; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_831 = 8'h3f == _t_T_2[23:16] ? 8'h75 : _GEN_830; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_832 = 8'h40 == _t_T_2[23:16] ? 8'h9 : _GEN_831; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_833 = 8'h41 == _t_T_2[23:16] ? 8'h83 : _GEN_832; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_834 = 8'h42 == _t_T_2[23:16] ? 8'h2c : _GEN_833; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_835 = 8'h43 == _t_T_2[23:16] ? 8'h1a : _GEN_834; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_836 = 8'h44 == _t_T_2[23:16] ? 8'h1b : _GEN_835; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_837 = 8'h45 == _t_T_2[23:16] ? 8'h6e : _GEN_836; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_838 = 8'h46 == _t_T_2[23:16] ? 8'h5a : _GEN_837; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_839 = 8'h47 == _t_T_2[23:16] ? 8'ha0 : _GEN_838; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_840 = 8'h48 == _t_T_2[23:16] ? 8'h52 : _GEN_839; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_841 = 8'h49 == _t_T_2[23:16] ? 8'h3b : _GEN_840; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_842 = 8'h4a == _t_T_2[23:16] ? 8'hd6 : _GEN_841; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_843 = 8'h4b == _t_T_2[23:16] ? 8'hb3 : _GEN_842; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_844 = 8'h4c == _t_T_2[23:16] ? 8'h29 : _GEN_843; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_845 = 8'h4d == _t_T_2[23:16] ? 8'he3 : _GEN_844; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_846 = 8'h4e == _t_T_2[23:16] ? 8'h2f : _GEN_845; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_847 = 8'h4f == _t_T_2[23:16] ? 8'h84 : _GEN_846; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_848 = 8'h50 == _t_T_2[23:16] ? 8'h53 : _GEN_847; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_849 = 8'h51 == _t_T_2[23:16] ? 8'hd1 : _GEN_848; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_850 = 8'h52 == _t_T_2[23:16] ? 8'h0 : _GEN_849; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_851 = 8'h53 == _t_T_2[23:16] ? 8'hed : _GEN_850; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_852 = 8'h54 == _t_T_2[23:16] ? 8'h20 : _GEN_851; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_853 = 8'h55 == _t_T_2[23:16] ? 8'hfc : _GEN_852; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_854 = 8'h56 == _t_T_2[23:16] ? 8'hb1 : _GEN_853; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_855 = 8'h57 == _t_T_2[23:16] ? 8'h5b : _GEN_854; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_856 = 8'h58 == _t_T_2[23:16] ? 8'h6a : _GEN_855; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_857 = 8'h59 == _t_T_2[23:16] ? 8'hcb : _GEN_856; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_858 = 8'h5a == _t_T_2[23:16] ? 8'hbe : _GEN_857; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_859 = 8'h5b == _t_T_2[23:16] ? 8'h39 : _GEN_858; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_860 = 8'h5c == _t_T_2[23:16] ? 8'h4a : _GEN_859; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_861 = 8'h5d == _t_T_2[23:16] ? 8'h4c : _GEN_860; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_862 = 8'h5e == _t_T_2[23:16] ? 8'h58 : _GEN_861; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_863 = 8'h5f == _t_T_2[23:16] ? 8'hcf : _GEN_862; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_864 = 8'h60 == _t_T_2[23:16] ? 8'hd0 : _GEN_863; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_865 = 8'h61 == _t_T_2[23:16] ? 8'hef : _GEN_864; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_866 = 8'h62 == _t_T_2[23:16] ? 8'haa : _GEN_865; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_867 = 8'h63 == _t_T_2[23:16] ? 8'hfb : _GEN_866; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_868 = 8'h64 == _t_T_2[23:16] ? 8'h43 : _GEN_867; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_869 = 8'h65 == _t_T_2[23:16] ? 8'h4d : _GEN_868; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_870 = 8'h66 == _t_T_2[23:16] ? 8'h33 : _GEN_869; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_871 = 8'h67 == _t_T_2[23:16] ? 8'h85 : _GEN_870; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_872 = 8'h68 == _t_T_2[23:16] ? 8'h45 : _GEN_871; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_873 = 8'h69 == _t_T_2[23:16] ? 8'hf9 : _GEN_872; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_874 = 8'h6a == _t_T_2[23:16] ? 8'h2 : _GEN_873; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_875 = 8'h6b == _t_T_2[23:16] ? 8'h7f : _GEN_874; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_876 = 8'h6c == _t_T_2[23:16] ? 8'h50 : _GEN_875; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_877 = 8'h6d == _t_T_2[23:16] ? 8'h3c : _GEN_876; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_878 = 8'h6e == _t_T_2[23:16] ? 8'h9f : _GEN_877; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_879 = 8'h6f == _t_T_2[23:16] ? 8'ha8 : _GEN_878; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_880 = 8'h70 == _t_T_2[23:16] ? 8'h51 : _GEN_879; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_881 = 8'h71 == _t_T_2[23:16] ? 8'ha3 : _GEN_880; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_882 = 8'h72 == _t_T_2[23:16] ? 8'h40 : _GEN_881; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_883 = 8'h73 == _t_T_2[23:16] ? 8'h8f : _GEN_882; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_884 = 8'h74 == _t_T_2[23:16] ? 8'h92 : _GEN_883; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_885 = 8'h75 == _t_T_2[23:16] ? 8'h9d : _GEN_884; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_886 = 8'h76 == _t_T_2[23:16] ? 8'h38 : _GEN_885; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_887 = 8'h77 == _t_T_2[23:16] ? 8'hf5 : _GEN_886; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_888 = 8'h78 == _t_T_2[23:16] ? 8'hbc : _GEN_887; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_889 = 8'h79 == _t_T_2[23:16] ? 8'hb6 : _GEN_888; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_890 = 8'h7a == _t_T_2[23:16] ? 8'hda : _GEN_889; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_891 = 8'h7b == _t_T_2[23:16] ? 8'h21 : _GEN_890; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_892 = 8'h7c == _t_T_2[23:16] ? 8'h10 : _GEN_891; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_893 = 8'h7d == _t_T_2[23:16] ? 8'hff : _GEN_892; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_894 = 8'h7e == _t_T_2[23:16] ? 8'hf3 : _GEN_893; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_895 = 8'h7f == _t_T_2[23:16] ? 8'hd2 : _GEN_894; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_896 = 8'h80 == _t_T_2[23:16] ? 8'hcd : _GEN_895; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_897 = 8'h81 == _t_T_2[23:16] ? 8'hc : _GEN_896; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_898 = 8'h82 == _t_T_2[23:16] ? 8'h13 : _GEN_897; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_899 = 8'h83 == _t_T_2[23:16] ? 8'hec : _GEN_898; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_900 = 8'h84 == _t_T_2[23:16] ? 8'h5f : _GEN_899; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_901 = 8'h85 == _t_T_2[23:16] ? 8'h97 : _GEN_900; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_902 = 8'h86 == _t_T_2[23:16] ? 8'h44 : _GEN_901; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_903 = 8'h87 == _t_T_2[23:16] ? 8'h17 : _GEN_902; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_904 = 8'h88 == _t_T_2[23:16] ? 8'hc4 : _GEN_903; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_905 = 8'h89 == _t_T_2[23:16] ? 8'ha7 : _GEN_904; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_906 = 8'h8a == _t_T_2[23:16] ? 8'h7e : _GEN_905; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_907 = 8'h8b == _t_T_2[23:16] ? 8'h3d : _GEN_906; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_908 = 8'h8c == _t_T_2[23:16] ? 8'h64 : _GEN_907; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_909 = 8'h8d == _t_T_2[23:16] ? 8'h5d : _GEN_908; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_910 = 8'h8e == _t_T_2[23:16] ? 8'h19 : _GEN_909; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_911 = 8'h8f == _t_T_2[23:16] ? 8'h73 : _GEN_910; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_912 = 8'h90 == _t_T_2[23:16] ? 8'h60 : _GEN_911; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_913 = 8'h91 == _t_T_2[23:16] ? 8'h81 : _GEN_912; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_914 = 8'h92 == _t_T_2[23:16] ? 8'h4f : _GEN_913; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_915 = 8'h93 == _t_T_2[23:16] ? 8'hdc : _GEN_914; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_916 = 8'h94 == _t_T_2[23:16] ? 8'h22 : _GEN_915; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_917 = 8'h95 == _t_T_2[23:16] ? 8'h2a : _GEN_916; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_918 = 8'h96 == _t_T_2[23:16] ? 8'h90 : _GEN_917; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_919 = 8'h97 == _t_T_2[23:16] ? 8'h88 : _GEN_918; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_920 = 8'h98 == _t_T_2[23:16] ? 8'h46 : _GEN_919; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_921 = 8'h99 == _t_T_2[23:16] ? 8'hee : _GEN_920; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_922 = 8'h9a == _t_T_2[23:16] ? 8'hb8 : _GEN_921; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_923 = 8'h9b == _t_T_2[23:16] ? 8'h14 : _GEN_922; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_924 = 8'h9c == _t_T_2[23:16] ? 8'hde : _GEN_923; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_925 = 8'h9d == _t_T_2[23:16] ? 8'h5e : _GEN_924; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_926 = 8'h9e == _t_T_2[23:16] ? 8'hb : _GEN_925; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_927 = 8'h9f == _t_T_2[23:16] ? 8'hdb : _GEN_926; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_928 = 8'ha0 == _t_T_2[23:16] ? 8'he0 : _GEN_927; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_929 = 8'ha1 == _t_T_2[23:16] ? 8'h32 : _GEN_928; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_930 = 8'ha2 == _t_T_2[23:16] ? 8'h3a : _GEN_929; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_931 = 8'ha3 == _t_T_2[23:16] ? 8'ha : _GEN_930; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_932 = 8'ha4 == _t_T_2[23:16] ? 8'h49 : _GEN_931; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_933 = 8'ha5 == _t_T_2[23:16] ? 8'h6 : _GEN_932; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_934 = 8'ha6 == _t_T_2[23:16] ? 8'h24 : _GEN_933; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_935 = 8'ha7 == _t_T_2[23:16] ? 8'h5c : _GEN_934; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_936 = 8'ha8 == _t_T_2[23:16] ? 8'hc2 : _GEN_935; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_937 = 8'ha9 == _t_T_2[23:16] ? 8'hd3 : _GEN_936; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_938 = 8'haa == _t_T_2[23:16] ? 8'hac : _GEN_937; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_939 = 8'hab == _t_T_2[23:16] ? 8'h62 : _GEN_938; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_940 = 8'hac == _t_T_2[23:16] ? 8'h91 : _GEN_939; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_941 = 8'had == _t_T_2[23:16] ? 8'h95 : _GEN_940; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_942 = 8'hae == _t_T_2[23:16] ? 8'he4 : _GEN_941; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_943 = 8'haf == _t_T_2[23:16] ? 8'h79 : _GEN_942; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_944 = 8'hb0 == _t_T_2[23:16] ? 8'he7 : _GEN_943; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_945 = 8'hb1 == _t_T_2[23:16] ? 8'hc8 : _GEN_944; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_946 = 8'hb2 == _t_T_2[23:16] ? 8'h37 : _GEN_945; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_947 = 8'hb3 == _t_T_2[23:16] ? 8'h6d : _GEN_946; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_948 = 8'hb4 == _t_T_2[23:16] ? 8'h8d : _GEN_947; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_949 = 8'hb5 == _t_T_2[23:16] ? 8'hd5 : _GEN_948; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_950 = 8'hb6 == _t_T_2[23:16] ? 8'h4e : _GEN_949; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_951 = 8'hb7 == _t_T_2[23:16] ? 8'ha9 : _GEN_950; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_952 = 8'hb8 == _t_T_2[23:16] ? 8'h6c : _GEN_951; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_953 = 8'hb9 == _t_T_2[23:16] ? 8'h56 : _GEN_952; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_954 = 8'hba == _t_T_2[23:16] ? 8'hf4 : _GEN_953; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_955 = 8'hbb == _t_T_2[23:16] ? 8'hea : _GEN_954; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_956 = 8'hbc == _t_T_2[23:16] ? 8'h65 : _GEN_955; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_957 = 8'hbd == _t_T_2[23:16] ? 8'h7a : _GEN_956; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_958 = 8'hbe == _t_T_2[23:16] ? 8'hae : _GEN_957; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_959 = 8'hbf == _t_T_2[23:16] ? 8'h8 : _GEN_958; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_960 = 8'hc0 == _t_T_2[23:16] ? 8'hba : _GEN_959; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_961 = 8'hc1 == _t_T_2[23:16] ? 8'h78 : _GEN_960; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_962 = 8'hc2 == _t_T_2[23:16] ? 8'h25 : _GEN_961; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_963 = 8'hc3 == _t_T_2[23:16] ? 8'h2e : _GEN_962; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_964 = 8'hc4 == _t_T_2[23:16] ? 8'h1c : _GEN_963; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_965 = 8'hc5 == _t_T_2[23:16] ? 8'ha6 : _GEN_964; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_966 = 8'hc6 == _t_T_2[23:16] ? 8'hb4 : _GEN_965; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_967 = 8'hc7 == _t_T_2[23:16] ? 8'hc6 : _GEN_966; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_968 = 8'hc8 == _t_T_2[23:16] ? 8'he8 : _GEN_967; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_969 = 8'hc9 == _t_T_2[23:16] ? 8'hdd : _GEN_968; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_970 = 8'hca == _t_T_2[23:16] ? 8'h74 : _GEN_969; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_971 = 8'hcb == _t_T_2[23:16] ? 8'h1f : _GEN_970; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_972 = 8'hcc == _t_T_2[23:16] ? 8'h4b : _GEN_971; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_973 = 8'hcd == _t_T_2[23:16] ? 8'hbd : _GEN_972; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_974 = 8'hce == _t_T_2[23:16] ? 8'h8b : _GEN_973; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_975 = 8'hcf == _t_T_2[23:16] ? 8'h8a : _GEN_974; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_976 = 8'hd0 == _t_T_2[23:16] ? 8'h70 : _GEN_975; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_977 = 8'hd1 == _t_T_2[23:16] ? 8'h3e : _GEN_976; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_978 = 8'hd2 == _t_T_2[23:16] ? 8'hb5 : _GEN_977; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_979 = 8'hd3 == _t_T_2[23:16] ? 8'h66 : _GEN_978; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_980 = 8'hd4 == _t_T_2[23:16] ? 8'h48 : _GEN_979; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_981 = 8'hd5 == _t_T_2[23:16] ? 8'h3 : _GEN_980; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_982 = 8'hd6 == _t_T_2[23:16] ? 8'hf6 : _GEN_981; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_983 = 8'hd7 == _t_T_2[23:16] ? 8'he : _GEN_982; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_984 = 8'hd8 == _t_T_2[23:16] ? 8'h61 : _GEN_983; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_985 = 8'hd9 == _t_T_2[23:16] ? 8'h35 : _GEN_984; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_986 = 8'hda == _t_T_2[23:16] ? 8'h57 : _GEN_985; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_987 = 8'hdb == _t_T_2[23:16] ? 8'hb9 : _GEN_986; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_988 = 8'hdc == _t_T_2[23:16] ? 8'h86 : _GEN_987; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_989 = 8'hdd == _t_T_2[23:16] ? 8'hc1 : _GEN_988; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_990 = 8'hde == _t_T_2[23:16] ? 8'h1d : _GEN_989; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_991 = 8'hdf == _t_T_2[23:16] ? 8'h9e : _GEN_990; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_992 = 8'he0 == _t_T_2[23:16] ? 8'he1 : _GEN_991; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_993 = 8'he1 == _t_T_2[23:16] ? 8'hf8 : _GEN_992; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_994 = 8'he2 == _t_T_2[23:16] ? 8'h98 : _GEN_993; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_995 = 8'he3 == _t_T_2[23:16] ? 8'h11 : _GEN_994; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_996 = 8'he4 == _t_T_2[23:16] ? 8'h69 : _GEN_995; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_997 = 8'he5 == _t_T_2[23:16] ? 8'hd9 : _GEN_996; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_998 = 8'he6 == _t_T_2[23:16] ? 8'h8e : _GEN_997; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_999 = 8'he7 == _t_T_2[23:16] ? 8'h94 : _GEN_998; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1000 = 8'he8 == _t_T_2[23:16] ? 8'h9b : _GEN_999; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1001 = 8'he9 == _t_T_2[23:16] ? 8'h1e : _GEN_1000; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1002 = 8'hea == _t_T_2[23:16] ? 8'h87 : _GEN_1001; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1003 = 8'heb == _t_T_2[23:16] ? 8'he9 : _GEN_1002; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1004 = 8'hec == _t_T_2[23:16] ? 8'hce : _GEN_1003; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1005 = 8'hed == _t_T_2[23:16] ? 8'h55 : _GEN_1004; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1006 = 8'hee == _t_T_2[23:16] ? 8'h28 : _GEN_1005; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1007 = 8'hef == _t_T_2[23:16] ? 8'hdf : _GEN_1006; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1008 = 8'hf0 == _t_T_2[23:16] ? 8'h8c : _GEN_1007; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1009 = 8'hf1 == _t_T_2[23:16] ? 8'ha1 : _GEN_1008; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1010 = 8'hf2 == _t_T_2[23:16] ? 8'h89 : _GEN_1009; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1011 = 8'hf3 == _t_T_2[23:16] ? 8'hd : _GEN_1010; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1012 = 8'hf4 == _t_T_2[23:16] ? 8'hbf : _GEN_1011; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1013 = 8'hf5 == _t_T_2[23:16] ? 8'he6 : _GEN_1012; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1014 = 8'hf6 == _t_T_2[23:16] ? 8'h42 : _GEN_1013; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1015 = 8'hf7 == _t_T_2[23:16] ? 8'h68 : _GEN_1014; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1016 = 8'hf8 == _t_T_2[23:16] ? 8'h41 : _GEN_1015; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1017 = 8'hf9 == _t_T_2[23:16] ? 8'h99 : _GEN_1016; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1018 = 8'hfa == _t_T_2[23:16] ? 8'h2d : _GEN_1017; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1019 = 8'hfb == _t_T_2[23:16] ? 8'hf : _GEN_1018; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1020 = 8'hfc == _t_T_2[23:16] ? 8'hb0 : _GEN_1019; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1021 = 8'hfd == _t_T_2[23:16] ? 8'h54 : _GEN_1020; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1022 = 8'hfe == _t_T_2[23:16] ? 8'hbb : _GEN_1021; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1023 = 8'hff == _t_T_2[23:16] ? 8'h16 : _GEN_1022; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [31:0] _t_T_7 = {_GEN_767,_GEN_1023,_GEN_255,_GEN_511}; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:8]
  wire [31:0] t = _t_T_7 ^ 32'h1000000; // @[src/main/scala/crypto/aes/KeySchedule.scala 59:32]
  wire [31:0] w_4 = w_0 ^ t; // @[src/main/scala/crypto/aes/KeySchedule.scala 63:21]
  wire [31:0] w_5 = w_1 ^ w_4; // @[src/main/scala/crypto/aes/KeySchedule.scala 63:21]
  wire [31:0] w_6 = w_2 ^ w_5; // @[src/main/scala/crypto/aes/KeySchedule.scala 63:21]
  wire [31:0] w_7 = w_3 ^ w_6; // @[src/main/scala/crypto/aes/KeySchedule.scala 63:21]
  wire [31:0] _t_T_10 = {w_7[23:0],w_7[31:24]}; // @[src/main/scala/crypto/aes/KeySchedule.scala 23:43]
  wire [7:0] _GEN_1025 = 8'h1 == _t_T_10[15:8] ? 8'h7c : 8'h63; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1026 = 8'h2 == _t_T_10[15:8] ? 8'h77 : _GEN_1025; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1027 = 8'h3 == _t_T_10[15:8] ? 8'h7b : _GEN_1026; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1028 = 8'h4 == _t_T_10[15:8] ? 8'hf2 : _GEN_1027; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1029 = 8'h5 == _t_T_10[15:8] ? 8'h6b : _GEN_1028; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1030 = 8'h6 == _t_T_10[15:8] ? 8'h6f : _GEN_1029; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1031 = 8'h7 == _t_T_10[15:8] ? 8'hc5 : _GEN_1030; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1032 = 8'h8 == _t_T_10[15:8] ? 8'h30 : _GEN_1031; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1033 = 8'h9 == _t_T_10[15:8] ? 8'h1 : _GEN_1032; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1034 = 8'ha == _t_T_10[15:8] ? 8'h67 : _GEN_1033; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1035 = 8'hb == _t_T_10[15:8] ? 8'h2b : _GEN_1034; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1036 = 8'hc == _t_T_10[15:8] ? 8'hfe : _GEN_1035; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1037 = 8'hd == _t_T_10[15:8] ? 8'hd7 : _GEN_1036; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1038 = 8'he == _t_T_10[15:8] ? 8'hab : _GEN_1037; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1039 = 8'hf == _t_T_10[15:8] ? 8'h76 : _GEN_1038; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1040 = 8'h10 == _t_T_10[15:8] ? 8'hca : _GEN_1039; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1041 = 8'h11 == _t_T_10[15:8] ? 8'h82 : _GEN_1040; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1042 = 8'h12 == _t_T_10[15:8] ? 8'hc9 : _GEN_1041; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1043 = 8'h13 == _t_T_10[15:8] ? 8'h7d : _GEN_1042; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1044 = 8'h14 == _t_T_10[15:8] ? 8'hfa : _GEN_1043; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1045 = 8'h15 == _t_T_10[15:8] ? 8'h59 : _GEN_1044; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1046 = 8'h16 == _t_T_10[15:8] ? 8'h47 : _GEN_1045; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1047 = 8'h17 == _t_T_10[15:8] ? 8'hf0 : _GEN_1046; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1048 = 8'h18 == _t_T_10[15:8] ? 8'had : _GEN_1047; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1049 = 8'h19 == _t_T_10[15:8] ? 8'hd4 : _GEN_1048; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1050 = 8'h1a == _t_T_10[15:8] ? 8'ha2 : _GEN_1049; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1051 = 8'h1b == _t_T_10[15:8] ? 8'haf : _GEN_1050; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1052 = 8'h1c == _t_T_10[15:8] ? 8'h9c : _GEN_1051; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1053 = 8'h1d == _t_T_10[15:8] ? 8'ha4 : _GEN_1052; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1054 = 8'h1e == _t_T_10[15:8] ? 8'h72 : _GEN_1053; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1055 = 8'h1f == _t_T_10[15:8] ? 8'hc0 : _GEN_1054; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1056 = 8'h20 == _t_T_10[15:8] ? 8'hb7 : _GEN_1055; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1057 = 8'h21 == _t_T_10[15:8] ? 8'hfd : _GEN_1056; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1058 = 8'h22 == _t_T_10[15:8] ? 8'h93 : _GEN_1057; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1059 = 8'h23 == _t_T_10[15:8] ? 8'h26 : _GEN_1058; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1060 = 8'h24 == _t_T_10[15:8] ? 8'h36 : _GEN_1059; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1061 = 8'h25 == _t_T_10[15:8] ? 8'h3f : _GEN_1060; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1062 = 8'h26 == _t_T_10[15:8] ? 8'hf7 : _GEN_1061; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1063 = 8'h27 == _t_T_10[15:8] ? 8'hcc : _GEN_1062; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1064 = 8'h28 == _t_T_10[15:8] ? 8'h34 : _GEN_1063; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1065 = 8'h29 == _t_T_10[15:8] ? 8'ha5 : _GEN_1064; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1066 = 8'h2a == _t_T_10[15:8] ? 8'he5 : _GEN_1065; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1067 = 8'h2b == _t_T_10[15:8] ? 8'hf1 : _GEN_1066; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1068 = 8'h2c == _t_T_10[15:8] ? 8'h71 : _GEN_1067; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1069 = 8'h2d == _t_T_10[15:8] ? 8'hd8 : _GEN_1068; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1070 = 8'h2e == _t_T_10[15:8] ? 8'h31 : _GEN_1069; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1071 = 8'h2f == _t_T_10[15:8] ? 8'h15 : _GEN_1070; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1072 = 8'h30 == _t_T_10[15:8] ? 8'h4 : _GEN_1071; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1073 = 8'h31 == _t_T_10[15:8] ? 8'hc7 : _GEN_1072; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1074 = 8'h32 == _t_T_10[15:8] ? 8'h23 : _GEN_1073; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1075 = 8'h33 == _t_T_10[15:8] ? 8'hc3 : _GEN_1074; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1076 = 8'h34 == _t_T_10[15:8] ? 8'h18 : _GEN_1075; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1077 = 8'h35 == _t_T_10[15:8] ? 8'h96 : _GEN_1076; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1078 = 8'h36 == _t_T_10[15:8] ? 8'h5 : _GEN_1077; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1079 = 8'h37 == _t_T_10[15:8] ? 8'h9a : _GEN_1078; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1080 = 8'h38 == _t_T_10[15:8] ? 8'h7 : _GEN_1079; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1081 = 8'h39 == _t_T_10[15:8] ? 8'h12 : _GEN_1080; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1082 = 8'h3a == _t_T_10[15:8] ? 8'h80 : _GEN_1081; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1083 = 8'h3b == _t_T_10[15:8] ? 8'he2 : _GEN_1082; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1084 = 8'h3c == _t_T_10[15:8] ? 8'heb : _GEN_1083; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1085 = 8'h3d == _t_T_10[15:8] ? 8'h27 : _GEN_1084; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1086 = 8'h3e == _t_T_10[15:8] ? 8'hb2 : _GEN_1085; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1087 = 8'h3f == _t_T_10[15:8] ? 8'h75 : _GEN_1086; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1088 = 8'h40 == _t_T_10[15:8] ? 8'h9 : _GEN_1087; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1089 = 8'h41 == _t_T_10[15:8] ? 8'h83 : _GEN_1088; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1090 = 8'h42 == _t_T_10[15:8] ? 8'h2c : _GEN_1089; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1091 = 8'h43 == _t_T_10[15:8] ? 8'h1a : _GEN_1090; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1092 = 8'h44 == _t_T_10[15:8] ? 8'h1b : _GEN_1091; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1093 = 8'h45 == _t_T_10[15:8] ? 8'h6e : _GEN_1092; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1094 = 8'h46 == _t_T_10[15:8] ? 8'h5a : _GEN_1093; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1095 = 8'h47 == _t_T_10[15:8] ? 8'ha0 : _GEN_1094; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1096 = 8'h48 == _t_T_10[15:8] ? 8'h52 : _GEN_1095; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1097 = 8'h49 == _t_T_10[15:8] ? 8'h3b : _GEN_1096; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1098 = 8'h4a == _t_T_10[15:8] ? 8'hd6 : _GEN_1097; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1099 = 8'h4b == _t_T_10[15:8] ? 8'hb3 : _GEN_1098; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1100 = 8'h4c == _t_T_10[15:8] ? 8'h29 : _GEN_1099; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1101 = 8'h4d == _t_T_10[15:8] ? 8'he3 : _GEN_1100; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1102 = 8'h4e == _t_T_10[15:8] ? 8'h2f : _GEN_1101; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1103 = 8'h4f == _t_T_10[15:8] ? 8'h84 : _GEN_1102; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1104 = 8'h50 == _t_T_10[15:8] ? 8'h53 : _GEN_1103; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1105 = 8'h51 == _t_T_10[15:8] ? 8'hd1 : _GEN_1104; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1106 = 8'h52 == _t_T_10[15:8] ? 8'h0 : _GEN_1105; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1107 = 8'h53 == _t_T_10[15:8] ? 8'hed : _GEN_1106; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1108 = 8'h54 == _t_T_10[15:8] ? 8'h20 : _GEN_1107; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1109 = 8'h55 == _t_T_10[15:8] ? 8'hfc : _GEN_1108; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1110 = 8'h56 == _t_T_10[15:8] ? 8'hb1 : _GEN_1109; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1111 = 8'h57 == _t_T_10[15:8] ? 8'h5b : _GEN_1110; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1112 = 8'h58 == _t_T_10[15:8] ? 8'h6a : _GEN_1111; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1113 = 8'h59 == _t_T_10[15:8] ? 8'hcb : _GEN_1112; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1114 = 8'h5a == _t_T_10[15:8] ? 8'hbe : _GEN_1113; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1115 = 8'h5b == _t_T_10[15:8] ? 8'h39 : _GEN_1114; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1116 = 8'h5c == _t_T_10[15:8] ? 8'h4a : _GEN_1115; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1117 = 8'h5d == _t_T_10[15:8] ? 8'h4c : _GEN_1116; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1118 = 8'h5e == _t_T_10[15:8] ? 8'h58 : _GEN_1117; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1119 = 8'h5f == _t_T_10[15:8] ? 8'hcf : _GEN_1118; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1120 = 8'h60 == _t_T_10[15:8] ? 8'hd0 : _GEN_1119; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1121 = 8'h61 == _t_T_10[15:8] ? 8'hef : _GEN_1120; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1122 = 8'h62 == _t_T_10[15:8] ? 8'haa : _GEN_1121; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1123 = 8'h63 == _t_T_10[15:8] ? 8'hfb : _GEN_1122; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1124 = 8'h64 == _t_T_10[15:8] ? 8'h43 : _GEN_1123; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1125 = 8'h65 == _t_T_10[15:8] ? 8'h4d : _GEN_1124; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1126 = 8'h66 == _t_T_10[15:8] ? 8'h33 : _GEN_1125; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1127 = 8'h67 == _t_T_10[15:8] ? 8'h85 : _GEN_1126; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1128 = 8'h68 == _t_T_10[15:8] ? 8'h45 : _GEN_1127; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1129 = 8'h69 == _t_T_10[15:8] ? 8'hf9 : _GEN_1128; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1130 = 8'h6a == _t_T_10[15:8] ? 8'h2 : _GEN_1129; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1131 = 8'h6b == _t_T_10[15:8] ? 8'h7f : _GEN_1130; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1132 = 8'h6c == _t_T_10[15:8] ? 8'h50 : _GEN_1131; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1133 = 8'h6d == _t_T_10[15:8] ? 8'h3c : _GEN_1132; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1134 = 8'h6e == _t_T_10[15:8] ? 8'h9f : _GEN_1133; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1135 = 8'h6f == _t_T_10[15:8] ? 8'ha8 : _GEN_1134; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1136 = 8'h70 == _t_T_10[15:8] ? 8'h51 : _GEN_1135; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1137 = 8'h71 == _t_T_10[15:8] ? 8'ha3 : _GEN_1136; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1138 = 8'h72 == _t_T_10[15:8] ? 8'h40 : _GEN_1137; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1139 = 8'h73 == _t_T_10[15:8] ? 8'h8f : _GEN_1138; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1140 = 8'h74 == _t_T_10[15:8] ? 8'h92 : _GEN_1139; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1141 = 8'h75 == _t_T_10[15:8] ? 8'h9d : _GEN_1140; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1142 = 8'h76 == _t_T_10[15:8] ? 8'h38 : _GEN_1141; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1143 = 8'h77 == _t_T_10[15:8] ? 8'hf5 : _GEN_1142; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1144 = 8'h78 == _t_T_10[15:8] ? 8'hbc : _GEN_1143; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1145 = 8'h79 == _t_T_10[15:8] ? 8'hb6 : _GEN_1144; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1146 = 8'h7a == _t_T_10[15:8] ? 8'hda : _GEN_1145; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1147 = 8'h7b == _t_T_10[15:8] ? 8'h21 : _GEN_1146; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1148 = 8'h7c == _t_T_10[15:8] ? 8'h10 : _GEN_1147; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1149 = 8'h7d == _t_T_10[15:8] ? 8'hff : _GEN_1148; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1150 = 8'h7e == _t_T_10[15:8] ? 8'hf3 : _GEN_1149; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1151 = 8'h7f == _t_T_10[15:8] ? 8'hd2 : _GEN_1150; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1152 = 8'h80 == _t_T_10[15:8] ? 8'hcd : _GEN_1151; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1153 = 8'h81 == _t_T_10[15:8] ? 8'hc : _GEN_1152; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1154 = 8'h82 == _t_T_10[15:8] ? 8'h13 : _GEN_1153; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1155 = 8'h83 == _t_T_10[15:8] ? 8'hec : _GEN_1154; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1156 = 8'h84 == _t_T_10[15:8] ? 8'h5f : _GEN_1155; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1157 = 8'h85 == _t_T_10[15:8] ? 8'h97 : _GEN_1156; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1158 = 8'h86 == _t_T_10[15:8] ? 8'h44 : _GEN_1157; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1159 = 8'h87 == _t_T_10[15:8] ? 8'h17 : _GEN_1158; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1160 = 8'h88 == _t_T_10[15:8] ? 8'hc4 : _GEN_1159; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1161 = 8'h89 == _t_T_10[15:8] ? 8'ha7 : _GEN_1160; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1162 = 8'h8a == _t_T_10[15:8] ? 8'h7e : _GEN_1161; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1163 = 8'h8b == _t_T_10[15:8] ? 8'h3d : _GEN_1162; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1164 = 8'h8c == _t_T_10[15:8] ? 8'h64 : _GEN_1163; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1165 = 8'h8d == _t_T_10[15:8] ? 8'h5d : _GEN_1164; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1166 = 8'h8e == _t_T_10[15:8] ? 8'h19 : _GEN_1165; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1167 = 8'h8f == _t_T_10[15:8] ? 8'h73 : _GEN_1166; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1168 = 8'h90 == _t_T_10[15:8] ? 8'h60 : _GEN_1167; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1169 = 8'h91 == _t_T_10[15:8] ? 8'h81 : _GEN_1168; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1170 = 8'h92 == _t_T_10[15:8] ? 8'h4f : _GEN_1169; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1171 = 8'h93 == _t_T_10[15:8] ? 8'hdc : _GEN_1170; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1172 = 8'h94 == _t_T_10[15:8] ? 8'h22 : _GEN_1171; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1173 = 8'h95 == _t_T_10[15:8] ? 8'h2a : _GEN_1172; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1174 = 8'h96 == _t_T_10[15:8] ? 8'h90 : _GEN_1173; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1175 = 8'h97 == _t_T_10[15:8] ? 8'h88 : _GEN_1174; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1176 = 8'h98 == _t_T_10[15:8] ? 8'h46 : _GEN_1175; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1177 = 8'h99 == _t_T_10[15:8] ? 8'hee : _GEN_1176; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1178 = 8'h9a == _t_T_10[15:8] ? 8'hb8 : _GEN_1177; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1179 = 8'h9b == _t_T_10[15:8] ? 8'h14 : _GEN_1178; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1180 = 8'h9c == _t_T_10[15:8] ? 8'hde : _GEN_1179; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1181 = 8'h9d == _t_T_10[15:8] ? 8'h5e : _GEN_1180; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1182 = 8'h9e == _t_T_10[15:8] ? 8'hb : _GEN_1181; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1183 = 8'h9f == _t_T_10[15:8] ? 8'hdb : _GEN_1182; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1184 = 8'ha0 == _t_T_10[15:8] ? 8'he0 : _GEN_1183; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1185 = 8'ha1 == _t_T_10[15:8] ? 8'h32 : _GEN_1184; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1186 = 8'ha2 == _t_T_10[15:8] ? 8'h3a : _GEN_1185; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1187 = 8'ha3 == _t_T_10[15:8] ? 8'ha : _GEN_1186; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1188 = 8'ha4 == _t_T_10[15:8] ? 8'h49 : _GEN_1187; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1189 = 8'ha5 == _t_T_10[15:8] ? 8'h6 : _GEN_1188; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1190 = 8'ha6 == _t_T_10[15:8] ? 8'h24 : _GEN_1189; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1191 = 8'ha7 == _t_T_10[15:8] ? 8'h5c : _GEN_1190; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1192 = 8'ha8 == _t_T_10[15:8] ? 8'hc2 : _GEN_1191; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1193 = 8'ha9 == _t_T_10[15:8] ? 8'hd3 : _GEN_1192; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1194 = 8'haa == _t_T_10[15:8] ? 8'hac : _GEN_1193; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1195 = 8'hab == _t_T_10[15:8] ? 8'h62 : _GEN_1194; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1196 = 8'hac == _t_T_10[15:8] ? 8'h91 : _GEN_1195; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1197 = 8'had == _t_T_10[15:8] ? 8'h95 : _GEN_1196; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1198 = 8'hae == _t_T_10[15:8] ? 8'he4 : _GEN_1197; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1199 = 8'haf == _t_T_10[15:8] ? 8'h79 : _GEN_1198; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1200 = 8'hb0 == _t_T_10[15:8] ? 8'he7 : _GEN_1199; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1201 = 8'hb1 == _t_T_10[15:8] ? 8'hc8 : _GEN_1200; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1202 = 8'hb2 == _t_T_10[15:8] ? 8'h37 : _GEN_1201; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1203 = 8'hb3 == _t_T_10[15:8] ? 8'h6d : _GEN_1202; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1204 = 8'hb4 == _t_T_10[15:8] ? 8'h8d : _GEN_1203; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1205 = 8'hb5 == _t_T_10[15:8] ? 8'hd5 : _GEN_1204; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1206 = 8'hb6 == _t_T_10[15:8] ? 8'h4e : _GEN_1205; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1207 = 8'hb7 == _t_T_10[15:8] ? 8'ha9 : _GEN_1206; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1208 = 8'hb8 == _t_T_10[15:8] ? 8'h6c : _GEN_1207; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1209 = 8'hb9 == _t_T_10[15:8] ? 8'h56 : _GEN_1208; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1210 = 8'hba == _t_T_10[15:8] ? 8'hf4 : _GEN_1209; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1211 = 8'hbb == _t_T_10[15:8] ? 8'hea : _GEN_1210; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1212 = 8'hbc == _t_T_10[15:8] ? 8'h65 : _GEN_1211; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1213 = 8'hbd == _t_T_10[15:8] ? 8'h7a : _GEN_1212; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1214 = 8'hbe == _t_T_10[15:8] ? 8'hae : _GEN_1213; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1215 = 8'hbf == _t_T_10[15:8] ? 8'h8 : _GEN_1214; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1216 = 8'hc0 == _t_T_10[15:8] ? 8'hba : _GEN_1215; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1217 = 8'hc1 == _t_T_10[15:8] ? 8'h78 : _GEN_1216; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1218 = 8'hc2 == _t_T_10[15:8] ? 8'h25 : _GEN_1217; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1219 = 8'hc3 == _t_T_10[15:8] ? 8'h2e : _GEN_1218; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1220 = 8'hc4 == _t_T_10[15:8] ? 8'h1c : _GEN_1219; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1221 = 8'hc5 == _t_T_10[15:8] ? 8'ha6 : _GEN_1220; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1222 = 8'hc6 == _t_T_10[15:8] ? 8'hb4 : _GEN_1221; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1223 = 8'hc7 == _t_T_10[15:8] ? 8'hc6 : _GEN_1222; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1224 = 8'hc8 == _t_T_10[15:8] ? 8'he8 : _GEN_1223; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1225 = 8'hc9 == _t_T_10[15:8] ? 8'hdd : _GEN_1224; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1226 = 8'hca == _t_T_10[15:8] ? 8'h74 : _GEN_1225; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1227 = 8'hcb == _t_T_10[15:8] ? 8'h1f : _GEN_1226; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1228 = 8'hcc == _t_T_10[15:8] ? 8'h4b : _GEN_1227; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1229 = 8'hcd == _t_T_10[15:8] ? 8'hbd : _GEN_1228; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1230 = 8'hce == _t_T_10[15:8] ? 8'h8b : _GEN_1229; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1231 = 8'hcf == _t_T_10[15:8] ? 8'h8a : _GEN_1230; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1232 = 8'hd0 == _t_T_10[15:8] ? 8'h70 : _GEN_1231; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1233 = 8'hd1 == _t_T_10[15:8] ? 8'h3e : _GEN_1232; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1234 = 8'hd2 == _t_T_10[15:8] ? 8'hb5 : _GEN_1233; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1235 = 8'hd3 == _t_T_10[15:8] ? 8'h66 : _GEN_1234; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1236 = 8'hd4 == _t_T_10[15:8] ? 8'h48 : _GEN_1235; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1237 = 8'hd5 == _t_T_10[15:8] ? 8'h3 : _GEN_1236; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1238 = 8'hd6 == _t_T_10[15:8] ? 8'hf6 : _GEN_1237; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1239 = 8'hd7 == _t_T_10[15:8] ? 8'he : _GEN_1238; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1240 = 8'hd8 == _t_T_10[15:8] ? 8'h61 : _GEN_1239; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1241 = 8'hd9 == _t_T_10[15:8] ? 8'h35 : _GEN_1240; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1242 = 8'hda == _t_T_10[15:8] ? 8'h57 : _GEN_1241; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1243 = 8'hdb == _t_T_10[15:8] ? 8'hb9 : _GEN_1242; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1244 = 8'hdc == _t_T_10[15:8] ? 8'h86 : _GEN_1243; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1245 = 8'hdd == _t_T_10[15:8] ? 8'hc1 : _GEN_1244; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1246 = 8'hde == _t_T_10[15:8] ? 8'h1d : _GEN_1245; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1247 = 8'hdf == _t_T_10[15:8] ? 8'h9e : _GEN_1246; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1248 = 8'he0 == _t_T_10[15:8] ? 8'he1 : _GEN_1247; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1249 = 8'he1 == _t_T_10[15:8] ? 8'hf8 : _GEN_1248; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1250 = 8'he2 == _t_T_10[15:8] ? 8'h98 : _GEN_1249; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1251 = 8'he3 == _t_T_10[15:8] ? 8'h11 : _GEN_1250; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1252 = 8'he4 == _t_T_10[15:8] ? 8'h69 : _GEN_1251; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1253 = 8'he5 == _t_T_10[15:8] ? 8'hd9 : _GEN_1252; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1254 = 8'he6 == _t_T_10[15:8] ? 8'h8e : _GEN_1253; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1255 = 8'he7 == _t_T_10[15:8] ? 8'h94 : _GEN_1254; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1256 = 8'he8 == _t_T_10[15:8] ? 8'h9b : _GEN_1255; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1257 = 8'he9 == _t_T_10[15:8] ? 8'h1e : _GEN_1256; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1258 = 8'hea == _t_T_10[15:8] ? 8'h87 : _GEN_1257; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1259 = 8'heb == _t_T_10[15:8] ? 8'he9 : _GEN_1258; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1260 = 8'hec == _t_T_10[15:8] ? 8'hce : _GEN_1259; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1261 = 8'hed == _t_T_10[15:8] ? 8'h55 : _GEN_1260; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1262 = 8'hee == _t_T_10[15:8] ? 8'h28 : _GEN_1261; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1263 = 8'hef == _t_T_10[15:8] ? 8'hdf : _GEN_1262; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1264 = 8'hf0 == _t_T_10[15:8] ? 8'h8c : _GEN_1263; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1265 = 8'hf1 == _t_T_10[15:8] ? 8'ha1 : _GEN_1264; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1266 = 8'hf2 == _t_T_10[15:8] ? 8'h89 : _GEN_1265; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1267 = 8'hf3 == _t_T_10[15:8] ? 8'hd : _GEN_1266; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1268 = 8'hf4 == _t_T_10[15:8] ? 8'hbf : _GEN_1267; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1269 = 8'hf5 == _t_T_10[15:8] ? 8'he6 : _GEN_1268; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1270 = 8'hf6 == _t_T_10[15:8] ? 8'h42 : _GEN_1269; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1271 = 8'hf7 == _t_T_10[15:8] ? 8'h68 : _GEN_1270; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1272 = 8'hf8 == _t_T_10[15:8] ? 8'h41 : _GEN_1271; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1273 = 8'hf9 == _t_T_10[15:8] ? 8'h99 : _GEN_1272; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1274 = 8'hfa == _t_T_10[15:8] ? 8'h2d : _GEN_1273; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1275 = 8'hfb == _t_T_10[15:8] ? 8'hf : _GEN_1274; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1276 = 8'hfc == _t_T_10[15:8] ? 8'hb0 : _GEN_1275; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1277 = 8'hfd == _t_T_10[15:8] ? 8'h54 : _GEN_1276; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1278 = 8'hfe == _t_T_10[15:8] ? 8'hbb : _GEN_1277; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1279 = 8'hff == _t_T_10[15:8] ? 8'h16 : _GEN_1278; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1281 = 8'h1 == _t_T_10[7:0] ? 8'h7c : 8'h63; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1282 = 8'h2 == _t_T_10[7:0] ? 8'h77 : _GEN_1281; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1283 = 8'h3 == _t_T_10[7:0] ? 8'h7b : _GEN_1282; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1284 = 8'h4 == _t_T_10[7:0] ? 8'hf2 : _GEN_1283; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1285 = 8'h5 == _t_T_10[7:0] ? 8'h6b : _GEN_1284; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1286 = 8'h6 == _t_T_10[7:0] ? 8'h6f : _GEN_1285; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1287 = 8'h7 == _t_T_10[7:0] ? 8'hc5 : _GEN_1286; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1288 = 8'h8 == _t_T_10[7:0] ? 8'h30 : _GEN_1287; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1289 = 8'h9 == _t_T_10[7:0] ? 8'h1 : _GEN_1288; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1290 = 8'ha == _t_T_10[7:0] ? 8'h67 : _GEN_1289; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1291 = 8'hb == _t_T_10[7:0] ? 8'h2b : _GEN_1290; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1292 = 8'hc == _t_T_10[7:0] ? 8'hfe : _GEN_1291; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1293 = 8'hd == _t_T_10[7:0] ? 8'hd7 : _GEN_1292; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1294 = 8'he == _t_T_10[7:0] ? 8'hab : _GEN_1293; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1295 = 8'hf == _t_T_10[7:0] ? 8'h76 : _GEN_1294; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1296 = 8'h10 == _t_T_10[7:0] ? 8'hca : _GEN_1295; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1297 = 8'h11 == _t_T_10[7:0] ? 8'h82 : _GEN_1296; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1298 = 8'h12 == _t_T_10[7:0] ? 8'hc9 : _GEN_1297; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1299 = 8'h13 == _t_T_10[7:0] ? 8'h7d : _GEN_1298; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1300 = 8'h14 == _t_T_10[7:0] ? 8'hfa : _GEN_1299; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1301 = 8'h15 == _t_T_10[7:0] ? 8'h59 : _GEN_1300; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1302 = 8'h16 == _t_T_10[7:0] ? 8'h47 : _GEN_1301; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1303 = 8'h17 == _t_T_10[7:0] ? 8'hf0 : _GEN_1302; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1304 = 8'h18 == _t_T_10[7:0] ? 8'had : _GEN_1303; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1305 = 8'h19 == _t_T_10[7:0] ? 8'hd4 : _GEN_1304; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1306 = 8'h1a == _t_T_10[7:0] ? 8'ha2 : _GEN_1305; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1307 = 8'h1b == _t_T_10[7:0] ? 8'haf : _GEN_1306; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1308 = 8'h1c == _t_T_10[7:0] ? 8'h9c : _GEN_1307; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1309 = 8'h1d == _t_T_10[7:0] ? 8'ha4 : _GEN_1308; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1310 = 8'h1e == _t_T_10[7:0] ? 8'h72 : _GEN_1309; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1311 = 8'h1f == _t_T_10[7:0] ? 8'hc0 : _GEN_1310; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1312 = 8'h20 == _t_T_10[7:0] ? 8'hb7 : _GEN_1311; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1313 = 8'h21 == _t_T_10[7:0] ? 8'hfd : _GEN_1312; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1314 = 8'h22 == _t_T_10[7:0] ? 8'h93 : _GEN_1313; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1315 = 8'h23 == _t_T_10[7:0] ? 8'h26 : _GEN_1314; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1316 = 8'h24 == _t_T_10[7:0] ? 8'h36 : _GEN_1315; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1317 = 8'h25 == _t_T_10[7:0] ? 8'h3f : _GEN_1316; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1318 = 8'h26 == _t_T_10[7:0] ? 8'hf7 : _GEN_1317; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1319 = 8'h27 == _t_T_10[7:0] ? 8'hcc : _GEN_1318; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1320 = 8'h28 == _t_T_10[7:0] ? 8'h34 : _GEN_1319; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1321 = 8'h29 == _t_T_10[7:0] ? 8'ha5 : _GEN_1320; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1322 = 8'h2a == _t_T_10[7:0] ? 8'he5 : _GEN_1321; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1323 = 8'h2b == _t_T_10[7:0] ? 8'hf1 : _GEN_1322; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1324 = 8'h2c == _t_T_10[7:0] ? 8'h71 : _GEN_1323; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1325 = 8'h2d == _t_T_10[7:0] ? 8'hd8 : _GEN_1324; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1326 = 8'h2e == _t_T_10[7:0] ? 8'h31 : _GEN_1325; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1327 = 8'h2f == _t_T_10[7:0] ? 8'h15 : _GEN_1326; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1328 = 8'h30 == _t_T_10[7:0] ? 8'h4 : _GEN_1327; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1329 = 8'h31 == _t_T_10[7:0] ? 8'hc7 : _GEN_1328; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1330 = 8'h32 == _t_T_10[7:0] ? 8'h23 : _GEN_1329; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1331 = 8'h33 == _t_T_10[7:0] ? 8'hc3 : _GEN_1330; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1332 = 8'h34 == _t_T_10[7:0] ? 8'h18 : _GEN_1331; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1333 = 8'h35 == _t_T_10[7:0] ? 8'h96 : _GEN_1332; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1334 = 8'h36 == _t_T_10[7:0] ? 8'h5 : _GEN_1333; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1335 = 8'h37 == _t_T_10[7:0] ? 8'h9a : _GEN_1334; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1336 = 8'h38 == _t_T_10[7:0] ? 8'h7 : _GEN_1335; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1337 = 8'h39 == _t_T_10[7:0] ? 8'h12 : _GEN_1336; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1338 = 8'h3a == _t_T_10[7:0] ? 8'h80 : _GEN_1337; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1339 = 8'h3b == _t_T_10[7:0] ? 8'he2 : _GEN_1338; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1340 = 8'h3c == _t_T_10[7:0] ? 8'heb : _GEN_1339; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1341 = 8'h3d == _t_T_10[7:0] ? 8'h27 : _GEN_1340; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1342 = 8'h3e == _t_T_10[7:0] ? 8'hb2 : _GEN_1341; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1343 = 8'h3f == _t_T_10[7:0] ? 8'h75 : _GEN_1342; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1344 = 8'h40 == _t_T_10[7:0] ? 8'h9 : _GEN_1343; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1345 = 8'h41 == _t_T_10[7:0] ? 8'h83 : _GEN_1344; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1346 = 8'h42 == _t_T_10[7:0] ? 8'h2c : _GEN_1345; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1347 = 8'h43 == _t_T_10[7:0] ? 8'h1a : _GEN_1346; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1348 = 8'h44 == _t_T_10[7:0] ? 8'h1b : _GEN_1347; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1349 = 8'h45 == _t_T_10[7:0] ? 8'h6e : _GEN_1348; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1350 = 8'h46 == _t_T_10[7:0] ? 8'h5a : _GEN_1349; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1351 = 8'h47 == _t_T_10[7:0] ? 8'ha0 : _GEN_1350; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1352 = 8'h48 == _t_T_10[7:0] ? 8'h52 : _GEN_1351; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1353 = 8'h49 == _t_T_10[7:0] ? 8'h3b : _GEN_1352; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1354 = 8'h4a == _t_T_10[7:0] ? 8'hd6 : _GEN_1353; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1355 = 8'h4b == _t_T_10[7:0] ? 8'hb3 : _GEN_1354; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1356 = 8'h4c == _t_T_10[7:0] ? 8'h29 : _GEN_1355; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1357 = 8'h4d == _t_T_10[7:0] ? 8'he3 : _GEN_1356; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1358 = 8'h4e == _t_T_10[7:0] ? 8'h2f : _GEN_1357; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1359 = 8'h4f == _t_T_10[7:0] ? 8'h84 : _GEN_1358; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1360 = 8'h50 == _t_T_10[7:0] ? 8'h53 : _GEN_1359; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1361 = 8'h51 == _t_T_10[7:0] ? 8'hd1 : _GEN_1360; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1362 = 8'h52 == _t_T_10[7:0] ? 8'h0 : _GEN_1361; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1363 = 8'h53 == _t_T_10[7:0] ? 8'hed : _GEN_1362; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1364 = 8'h54 == _t_T_10[7:0] ? 8'h20 : _GEN_1363; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1365 = 8'h55 == _t_T_10[7:0] ? 8'hfc : _GEN_1364; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1366 = 8'h56 == _t_T_10[7:0] ? 8'hb1 : _GEN_1365; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1367 = 8'h57 == _t_T_10[7:0] ? 8'h5b : _GEN_1366; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1368 = 8'h58 == _t_T_10[7:0] ? 8'h6a : _GEN_1367; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1369 = 8'h59 == _t_T_10[7:0] ? 8'hcb : _GEN_1368; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1370 = 8'h5a == _t_T_10[7:0] ? 8'hbe : _GEN_1369; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1371 = 8'h5b == _t_T_10[7:0] ? 8'h39 : _GEN_1370; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1372 = 8'h5c == _t_T_10[7:0] ? 8'h4a : _GEN_1371; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1373 = 8'h5d == _t_T_10[7:0] ? 8'h4c : _GEN_1372; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1374 = 8'h5e == _t_T_10[7:0] ? 8'h58 : _GEN_1373; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1375 = 8'h5f == _t_T_10[7:0] ? 8'hcf : _GEN_1374; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1376 = 8'h60 == _t_T_10[7:0] ? 8'hd0 : _GEN_1375; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1377 = 8'h61 == _t_T_10[7:0] ? 8'hef : _GEN_1376; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1378 = 8'h62 == _t_T_10[7:0] ? 8'haa : _GEN_1377; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1379 = 8'h63 == _t_T_10[7:0] ? 8'hfb : _GEN_1378; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1380 = 8'h64 == _t_T_10[7:0] ? 8'h43 : _GEN_1379; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1381 = 8'h65 == _t_T_10[7:0] ? 8'h4d : _GEN_1380; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1382 = 8'h66 == _t_T_10[7:0] ? 8'h33 : _GEN_1381; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1383 = 8'h67 == _t_T_10[7:0] ? 8'h85 : _GEN_1382; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1384 = 8'h68 == _t_T_10[7:0] ? 8'h45 : _GEN_1383; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1385 = 8'h69 == _t_T_10[7:0] ? 8'hf9 : _GEN_1384; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1386 = 8'h6a == _t_T_10[7:0] ? 8'h2 : _GEN_1385; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1387 = 8'h6b == _t_T_10[7:0] ? 8'h7f : _GEN_1386; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1388 = 8'h6c == _t_T_10[7:0] ? 8'h50 : _GEN_1387; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1389 = 8'h6d == _t_T_10[7:0] ? 8'h3c : _GEN_1388; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1390 = 8'h6e == _t_T_10[7:0] ? 8'h9f : _GEN_1389; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1391 = 8'h6f == _t_T_10[7:0] ? 8'ha8 : _GEN_1390; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1392 = 8'h70 == _t_T_10[7:0] ? 8'h51 : _GEN_1391; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1393 = 8'h71 == _t_T_10[7:0] ? 8'ha3 : _GEN_1392; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1394 = 8'h72 == _t_T_10[7:0] ? 8'h40 : _GEN_1393; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1395 = 8'h73 == _t_T_10[7:0] ? 8'h8f : _GEN_1394; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1396 = 8'h74 == _t_T_10[7:0] ? 8'h92 : _GEN_1395; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1397 = 8'h75 == _t_T_10[7:0] ? 8'h9d : _GEN_1396; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1398 = 8'h76 == _t_T_10[7:0] ? 8'h38 : _GEN_1397; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1399 = 8'h77 == _t_T_10[7:0] ? 8'hf5 : _GEN_1398; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1400 = 8'h78 == _t_T_10[7:0] ? 8'hbc : _GEN_1399; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1401 = 8'h79 == _t_T_10[7:0] ? 8'hb6 : _GEN_1400; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1402 = 8'h7a == _t_T_10[7:0] ? 8'hda : _GEN_1401; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1403 = 8'h7b == _t_T_10[7:0] ? 8'h21 : _GEN_1402; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1404 = 8'h7c == _t_T_10[7:0] ? 8'h10 : _GEN_1403; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1405 = 8'h7d == _t_T_10[7:0] ? 8'hff : _GEN_1404; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1406 = 8'h7e == _t_T_10[7:0] ? 8'hf3 : _GEN_1405; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1407 = 8'h7f == _t_T_10[7:0] ? 8'hd2 : _GEN_1406; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1408 = 8'h80 == _t_T_10[7:0] ? 8'hcd : _GEN_1407; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1409 = 8'h81 == _t_T_10[7:0] ? 8'hc : _GEN_1408; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1410 = 8'h82 == _t_T_10[7:0] ? 8'h13 : _GEN_1409; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1411 = 8'h83 == _t_T_10[7:0] ? 8'hec : _GEN_1410; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1412 = 8'h84 == _t_T_10[7:0] ? 8'h5f : _GEN_1411; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1413 = 8'h85 == _t_T_10[7:0] ? 8'h97 : _GEN_1412; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1414 = 8'h86 == _t_T_10[7:0] ? 8'h44 : _GEN_1413; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1415 = 8'h87 == _t_T_10[7:0] ? 8'h17 : _GEN_1414; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1416 = 8'h88 == _t_T_10[7:0] ? 8'hc4 : _GEN_1415; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1417 = 8'h89 == _t_T_10[7:0] ? 8'ha7 : _GEN_1416; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1418 = 8'h8a == _t_T_10[7:0] ? 8'h7e : _GEN_1417; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1419 = 8'h8b == _t_T_10[7:0] ? 8'h3d : _GEN_1418; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1420 = 8'h8c == _t_T_10[7:0] ? 8'h64 : _GEN_1419; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1421 = 8'h8d == _t_T_10[7:0] ? 8'h5d : _GEN_1420; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1422 = 8'h8e == _t_T_10[7:0] ? 8'h19 : _GEN_1421; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1423 = 8'h8f == _t_T_10[7:0] ? 8'h73 : _GEN_1422; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1424 = 8'h90 == _t_T_10[7:0] ? 8'h60 : _GEN_1423; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1425 = 8'h91 == _t_T_10[7:0] ? 8'h81 : _GEN_1424; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1426 = 8'h92 == _t_T_10[7:0] ? 8'h4f : _GEN_1425; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1427 = 8'h93 == _t_T_10[7:0] ? 8'hdc : _GEN_1426; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1428 = 8'h94 == _t_T_10[7:0] ? 8'h22 : _GEN_1427; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1429 = 8'h95 == _t_T_10[7:0] ? 8'h2a : _GEN_1428; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1430 = 8'h96 == _t_T_10[7:0] ? 8'h90 : _GEN_1429; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1431 = 8'h97 == _t_T_10[7:0] ? 8'h88 : _GEN_1430; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1432 = 8'h98 == _t_T_10[7:0] ? 8'h46 : _GEN_1431; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1433 = 8'h99 == _t_T_10[7:0] ? 8'hee : _GEN_1432; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1434 = 8'h9a == _t_T_10[7:0] ? 8'hb8 : _GEN_1433; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1435 = 8'h9b == _t_T_10[7:0] ? 8'h14 : _GEN_1434; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1436 = 8'h9c == _t_T_10[7:0] ? 8'hde : _GEN_1435; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1437 = 8'h9d == _t_T_10[7:0] ? 8'h5e : _GEN_1436; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1438 = 8'h9e == _t_T_10[7:0] ? 8'hb : _GEN_1437; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1439 = 8'h9f == _t_T_10[7:0] ? 8'hdb : _GEN_1438; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1440 = 8'ha0 == _t_T_10[7:0] ? 8'he0 : _GEN_1439; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1441 = 8'ha1 == _t_T_10[7:0] ? 8'h32 : _GEN_1440; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1442 = 8'ha2 == _t_T_10[7:0] ? 8'h3a : _GEN_1441; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1443 = 8'ha3 == _t_T_10[7:0] ? 8'ha : _GEN_1442; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1444 = 8'ha4 == _t_T_10[7:0] ? 8'h49 : _GEN_1443; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1445 = 8'ha5 == _t_T_10[7:0] ? 8'h6 : _GEN_1444; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1446 = 8'ha6 == _t_T_10[7:0] ? 8'h24 : _GEN_1445; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1447 = 8'ha7 == _t_T_10[7:0] ? 8'h5c : _GEN_1446; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1448 = 8'ha8 == _t_T_10[7:0] ? 8'hc2 : _GEN_1447; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1449 = 8'ha9 == _t_T_10[7:0] ? 8'hd3 : _GEN_1448; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1450 = 8'haa == _t_T_10[7:0] ? 8'hac : _GEN_1449; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1451 = 8'hab == _t_T_10[7:0] ? 8'h62 : _GEN_1450; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1452 = 8'hac == _t_T_10[7:0] ? 8'h91 : _GEN_1451; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1453 = 8'had == _t_T_10[7:0] ? 8'h95 : _GEN_1452; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1454 = 8'hae == _t_T_10[7:0] ? 8'he4 : _GEN_1453; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1455 = 8'haf == _t_T_10[7:0] ? 8'h79 : _GEN_1454; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1456 = 8'hb0 == _t_T_10[7:0] ? 8'he7 : _GEN_1455; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1457 = 8'hb1 == _t_T_10[7:0] ? 8'hc8 : _GEN_1456; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1458 = 8'hb2 == _t_T_10[7:0] ? 8'h37 : _GEN_1457; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1459 = 8'hb3 == _t_T_10[7:0] ? 8'h6d : _GEN_1458; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1460 = 8'hb4 == _t_T_10[7:0] ? 8'h8d : _GEN_1459; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1461 = 8'hb5 == _t_T_10[7:0] ? 8'hd5 : _GEN_1460; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1462 = 8'hb6 == _t_T_10[7:0] ? 8'h4e : _GEN_1461; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1463 = 8'hb7 == _t_T_10[7:0] ? 8'ha9 : _GEN_1462; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1464 = 8'hb8 == _t_T_10[7:0] ? 8'h6c : _GEN_1463; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1465 = 8'hb9 == _t_T_10[7:0] ? 8'h56 : _GEN_1464; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1466 = 8'hba == _t_T_10[7:0] ? 8'hf4 : _GEN_1465; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1467 = 8'hbb == _t_T_10[7:0] ? 8'hea : _GEN_1466; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1468 = 8'hbc == _t_T_10[7:0] ? 8'h65 : _GEN_1467; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1469 = 8'hbd == _t_T_10[7:0] ? 8'h7a : _GEN_1468; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1470 = 8'hbe == _t_T_10[7:0] ? 8'hae : _GEN_1469; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1471 = 8'hbf == _t_T_10[7:0] ? 8'h8 : _GEN_1470; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1472 = 8'hc0 == _t_T_10[7:0] ? 8'hba : _GEN_1471; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1473 = 8'hc1 == _t_T_10[7:0] ? 8'h78 : _GEN_1472; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1474 = 8'hc2 == _t_T_10[7:0] ? 8'h25 : _GEN_1473; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1475 = 8'hc3 == _t_T_10[7:0] ? 8'h2e : _GEN_1474; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1476 = 8'hc4 == _t_T_10[7:0] ? 8'h1c : _GEN_1475; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1477 = 8'hc5 == _t_T_10[7:0] ? 8'ha6 : _GEN_1476; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1478 = 8'hc6 == _t_T_10[7:0] ? 8'hb4 : _GEN_1477; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1479 = 8'hc7 == _t_T_10[7:0] ? 8'hc6 : _GEN_1478; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1480 = 8'hc8 == _t_T_10[7:0] ? 8'he8 : _GEN_1479; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1481 = 8'hc9 == _t_T_10[7:0] ? 8'hdd : _GEN_1480; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1482 = 8'hca == _t_T_10[7:0] ? 8'h74 : _GEN_1481; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1483 = 8'hcb == _t_T_10[7:0] ? 8'h1f : _GEN_1482; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1484 = 8'hcc == _t_T_10[7:0] ? 8'h4b : _GEN_1483; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1485 = 8'hcd == _t_T_10[7:0] ? 8'hbd : _GEN_1484; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1486 = 8'hce == _t_T_10[7:0] ? 8'h8b : _GEN_1485; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1487 = 8'hcf == _t_T_10[7:0] ? 8'h8a : _GEN_1486; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1488 = 8'hd0 == _t_T_10[7:0] ? 8'h70 : _GEN_1487; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1489 = 8'hd1 == _t_T_10[7:0] ? 8'h3e : _GEN_1488; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1490 = 8'hd2 == _t_T_10[7:0] ? 8'hb5 : _GEN_1489; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1491 = 8'hd3 == _t_T_10[7:0] ? 8'h66 : _GEN_1490; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1492 = 8'hd4 == _t_T_10[7:0] ? 8'h48 : _GEN_1491; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1493 = 8'hd5 == _t_T_10[7:0] ? 8'h3 : _GEN_1492; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1494 = 8'hd6 == _t_T_10[7:0] ? 8'hf6 : _GEN_1493; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1495 = 8'hd7 == _t_T_10[7:0] ? 8'he : _GEN_1494; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1496 = 8'hd8 == _t_T_10[7:0] ? 8'h61 : _GEN_1495; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1497 = 8'hd9 == _t_T_10[7:0] ? 8'h35 : _GEN_1496; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1498 = 8'hda == _t_T_10[7:0] ? 8'h57 : _GEN_1497; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1499 = 8'hdb == _t_T_10[7:0] ? 8'hb9 : _GEN_1498; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1500 = 8'hdc == _t_T_10[7:0] ? 8'h86 : _GEN_1499; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1501 = 8'hdd == _t_T_10[7:0] ? 8'hc1 : _GEN_1500; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1502 = 8'hde == _t_T_10[7:0] ? 8'h1d : _GEN_1501; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1503 = 8'hdf == _t_T_10[7:0] ? 8'h9e : _GEN_1502; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1504 = 8'he0 == _t_T_10[7:0] ? 8'he1 : _GEN_1503; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1505 = 8'he1 == _t_T_10[7:0] ? 8'hf8 : _GEN_1504; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1506 = 8'he2 == _t_T_10[7:0] ? 8'h98 : _GEN_1505; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1507 = 8'he3 == _t_T_10[7:0] ? 8'h11 : _GEN_1506; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1508 = 8'he4 == _t_T_10[7:0] ? 8'h69 : _GEN_1507; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1509 = 8'he5 == _t_T_10[7:0] ? 8'hd9 : _GEN_1508; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1510 = 8'he6 == _t_T_10[7:0] ? 8'h8e : _GEN_1509; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1511 = 8'he7 == _t_T_10[7:0] ? 8'h94 : _GEN_1510; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1512 = 8'he8 == _t_T_10[7:0] ? 8'h9b : _GEN_1511; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1513 = 8'he9 == _t_T_10[7:0] ? 8'h1e : _GEN_1512; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1514 = 8'hea == _t_T_10[7:0] ? 8'h87 : _GEN_1513; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1515 = 8'heb == _t_T_10[7:0] ? 8'he9 : _GEN_1514; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1516 = 8'hec == _t_T_10[7:0] ? 8'hce : _GEN_1515; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1517 = 8'hed == _t_T_10[7:0] ? 8'h55 : _GEN_1516; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1518 = 8'hee == _t_T_10[7:0] ? 8'h28 : _GEN_1517; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1519 = 8'hef == _t_T_10[7:0] ? 8'hdf : _GEN_1518; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1520 = 8'hf0 == _t_T_10[7:0] ? 8'h8c : _GEN_1519; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1521 = 8'hf1 == _t_T_10[7:0] ? 8'ha1 : _GEN_1520; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1522 = 8'hf2 == _t_T_10[7:0] ? 8'h89 : _GEN_1521; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1523 = 8'hf3 == _t_T_10[7:0] ? 8'hd : _GEN_1522; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1524 = 8'hf4 == _t_T_10[7:0] ? 8'hbf : _GEN_1523; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1525 = 8'hf5 == _t_T_10[7:0] ? 8'he6 : _GEN_1524; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1526 = 8'hf6 == _t_T_10[7:0] ? 8'h42 : _GEN_1525; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1527 = 8'hf7 == _t_T_10[7:0] ? 8'h68 : _GEN_1526; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1528 = 8'hf8 == _t_T_10[7:0] ? 8'h41 : _GEN_1527; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1529 = 8'hf9 == _t_T_10[7:0] ? 8'h99 : _GEN_1528; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1530 = 8'hfa == _t_T_10[7:0] ? 8'h2d : _GEN_1529; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1531 = 8'hfb == _t_T_10[7:0] ? 8'hf : _GEN_1530; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1532 = 8'hfc == _t_T_10[7:0] ? 8'hb0 : _GEN_1531; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1533 = 8'hfd == _t_T_10[7:0] ? 8'h54 : _GEN_1532; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1534 = 8'hfe == _t_T_10[7:0] ? 8'hbb : _GEN_1533; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1535 = 8'hff == _t_T_10[7:0] ? 8'h16 : _GEN_1534; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1537 = 8'h1 == _t_T_10[31:24] ? 8'h7c : 8'h63; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1538 = 8'h2 == _t_T_10[31:24] ? 8'h77 : _GEN_1537; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1539 = 8'h3 == _t_T_10[31:24] ? 8'h7b : _GEN_1538; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1540 = 8'h4 == _t_T_10[31:24] ? 8'hf2 : _GEN_1539; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1541 = 8'h5 == _t_T_10[31:24] ? 8'h6b : _GEN_1540; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1542 = 8'h6 == _t_T_10[31:24] ? 8'h6f : _GEN_1541; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1543 = 8'h7 == _t_T_10[31:24] ? 8'hc5 : _GEN_1542; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1544 = 8'h8 == _t_T_10[31:24] ? 8'h30 : _GEN_1543; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1545 = 8'h9 == _t_T_10[31:24] ? 8'h1 : _GEN_1544; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1546 = 8'ha == _t_T_10[31:24] ? 8'h67 : _GEN_1545; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1547 = 8'hb == _t_T_10[31:24] ? 8'h2b : _GEN_1546; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1548 = 8'hc == _t_T_10[31:24] ? 8'hfe : _GEN_1547; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1549 = 8'hd == _t_T_10[31:24] ? 8'hd7 : _GEN_1548; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1550 = 8'he == _t_T_10[31:24] ? 8'hab : _GEN_1549; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1551 = 8'hf == _t_T_10[31:24] ? 8'h76 : _GEN_1550; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1552 = 8'h10 == _t_T_10[31:24] ? 8'hca : _GEN_1551; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1553 = 8'h11 == _t_T_10[31:24] ? 8'h82 : _GEN_1552; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1554 = 8'h12 == _t_T_10[31:24] ? 8'hc9 : _GEN_1553; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1555 = 8'h13 == _t_T_10[31:24] ? 8'h7d : _GEN_1554; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1556 = 8'h14 == _t_T_10[31:24] ? 8'hfa : _GEN_1555; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1557 = 8'h15 == _t_T_10[31:24] ? 8'h59 : _GEN_1556; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1558 = 8'h16 == _t_T_10[31:24] ? 8'h47 : _GEN_1557; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1559 = 8'h17 == _t_T_10[31:24] ? 8'hf0 : _GEN_1558; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1560 = 8'h18 == _t_T_10[31:24] ? 8'had : _GEN_1559; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1561 = 8'h19 == _t_T_10[31:24] ? 8'hd4 : _GEN_1560; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1562 = 8'h1a == _t_T_10[31:24] ? 8'ha2 : _GEN_1561; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1563 = 8'h1b == _t_T_10[31:24] ? 8'haf : _GEN_1562; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1564 = 8'h1c == _t_T_10[31:24] ? 8'h9c : _GEN_1563; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1565 = 8'h1d == _t_T_10[31:24] ? 8'ha4 : _GEN_1564; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1566 = 8'h1e == _t_T_10[31:24] ? 8'h72 : _GEN_1565; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1567 = 8'h1f == _t_T_10[31:24] ? 8'hc0 : _GEN_1566; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1568 = 8'h20 == _t_T_10[31:24] ? 8'hb7 : _GEN_1567; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1569 = 8'h21 == _t_T_10[31:24] ? 8'hfd : _GEN_1568; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1570 = 8'h22 == _t_T_10[31:24] ? 8'h93 : _GEN_1569; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1571 = 8'h23 == _t_T_10[31:24] ? 8'h26 : _GEN_1570; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1572 = 8'h24 == _t_T_10[31:24] ? 8'h36 : _GEN_1571; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1573 = 8'h25 == _t_T_10[31:24] ? 8'h3f : _GEN_1572; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1574 = 8'h26 == _t_T_10[31:24] ? 8'hf7 : _GEN_1573; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1575 = 8'h27 == _t_T_10[31:24] ? 8'hcc : _GEN_1574; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1576 = 8'h28 == _t_T_10[31:24] ? 8'h34 : _GEN_1575; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1577 = 8'h29 == _t_T_10[31:24] ? 8'ha5 : _GEN_1576; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1578 = 8'h2a == _t_T_10[31:24] ? 8'he5 : _GEN_1577; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1579 = 8'h2b == _t_T_10[31:24] ? 8'hf1 : _GEN_1578; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1580 = 8'h2c == _t_T_10[31:24] ? 8'h71 : _GEN_1579; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1581 = 8'h2d == _t_T_10[31:24] ? 8'hd8 : _GEN_1580; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1582 = 8'h2e == _t_T_10[31:24] ? 8'h31 : _GEN_1581; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1583 = 8'h2f == _t_T_10[31:24] ? 8'h15 : _GEN_1582; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1584 = 8'h30 == _t_T_10[31:24] ? 8'h4 : _GEN_1583; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1585 = 8'h31 == _t_T_10[31:24] ? 8'hc7 : _GEN_1584; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1586 = 8'h32 == _t_T_10[31:24] ? 8'h23 : _GEN_1585; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1587 = 8'h33 == _t_T_10[31:24] ? 8'hc3 : _GEN_1586; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1588 = 8'h34 == _t_T_10[31:24] ? 8'h18 : _GEN_1587; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1589 = 8'h35 == _t_T_10[31:24] ? 8'h96 : _GEN_1588; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1590 = 8'h36 == _t_T_10[31:24] ? 8'h5 : _GEN_1589; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1591 = 8'h37 == _t_T_10[31:24] ? 8'h9a : _GEN_1590; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1592 = 8'h38 == _t_T_10[31:24] ? 8'h7 : _GEN_1591; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1593 = 8'h39 == _t_T_10[31:24] ? 8'h12 : _GEN_1592; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1594 = 8'h3a == _t_T_10[31:24] ? 8'h80 : _GEN_1593; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1595 = 8'h3b == _t_T_10[31:24] ? 8'he2 : _GEN_1594; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1596 = 8'h3c == _t_T_10[31:24] ? 8'heb : _GEN_1595; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1597 = 8'h3d == _t_T_10[31:24] ? 8'h27 : _GEN_1596; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1598 = 8'h3e == _t_T_10[31:24] ? 8'hb2 : _GEN_1597; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1599 = 8'h3f == _t_T_10[31:24] ? 8'h75 : _GEN_1598; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1600 = 8'h40 == _t_T_10[31:24] ? 8'h9 : _GEN_1599; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1601 = 8'h41 == _t_T_10[31:24] ? 8'h83 : _GEN_1600; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1602 = 8'h42 == _t_T_10[31:24] ? 8'h2c : _GEN_1601; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1603 = 8'h43 == _t_T_10[31:24] ? 8'h1a : _GEN_1602; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1604 = 8'h44 == _t_T_10[31:24] ? 8'h1b : _GEN_1603; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1605 = 8'h45 == _t_T_10[31:24] ? 8'h6e : _GEN_1604; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1606 = 8'h46 == _t_T_10[31:24] ? 8'h5a : _GEN_1605; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1607 = 8'h47 == _t_T_10[31:24] ? 8'ha0 : _GEN_1606; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1608 = 8'h48 == _t_T_10[31:24] ? 8'h52 : _GEN_1607; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1609 = 8'h49 == _t_T_10[31:24] ? 8'h3b : _GEN_1608; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1610 = 8'h4a == _t_T_10[31:24] ? 8'hd6 : _GEN_1609; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1611 = 8'h4b == _t_T_10[31:24] ? 8'hb3 : _GEN_1610; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1612 = 8'h4c == _t_T_10[31:24] ? 8'h29 : _GEN_1611; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1613 = 8'h4d == _t_T_10[31:24] ? 8'he3 : _GEN_1612; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1614 = 8'h4e == _t_T_10[31:24] ? 8'h2f : _GEN_1613; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1615 = 8'h4f == _t_T_10[31:24] ? 8'h84 : _GEN_1614; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1616 = 8'h50 == _t_T_10[31:24] ? 8'h53 : _GEN_1615; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1617 = 8'h51 == _t_T_10[31:24] ? 8'hd1 : _GEN_1616; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1618 = 8'h52 == _t_T_10[31:24] ? 8'h0 : _GEN_1617; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1619 = 8'h53 == _t_T_10[31:24] ? 8'hed : _GEN_1618; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1620 = 8'h54 == _t_T_10[31:24] ? 8'h20 : _GEN_1619; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1621 = 8'h55 == _t_T_10[31:24] ? 8'hfc : _GEN_1620; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1622 = 8'h56 == _t_T_10[31:24] ? 8'hb1 : _GEN_1621; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1623 = 8'h57 == _t_T_10[31:24] ? 8'h5b : _GEN_1622; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1624 = 8'h58 == _t_T_10[31:24] ? 8'h6a : _GEN_1623; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1625 = 8'h59 == _t_T_10[31:24] ? 8'hcb : _GEN_1624; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1626 = 8'h5a == _t_T_10[31:24] ? 8'hbe : _GEN_1625; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1627 = 8'h5b == _t_T_10[31:24] ? 8'h39 : _GEN_1626; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1628 = 8'h5c == _t_T_10[31:24] ? 8'h4a : _GEN_1627; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1629 = 8'h5d == _t_T_10[31:24] ? 8'h4c : _GEN_1628; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1630 = 8'h5e == _t_T_10[31:24] ? 8'h58 : _GEN_1629; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1631 = 8'h5f == _t_T_10[31:24] ? 8'hcf : _GEN_1630; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1632 = 8'h60 == _t_T_10[31:24] ? 8'hd0 : _GEN_1631; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1633 = 8'h61 == _t_T_10[31:24] ? 8'hef : _GEN_1632; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1634 = 8'h62 == _t_T_10[31:24] ? 8'haa : _GEN_1633; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1635 = 8'h63 == _t_T_10[31:24] ? 8'hfb : _GEN_1634; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1636 = 8'h64 == _t_T_10[31:24] ? 8'h43 : _GEN_1635; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1637 = 8'h65 == _t_T_10[31:24] ? 8'h4d : _GEN_1636; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1638 = 8'h66 == _t_T_10[31:24] ? 8'h33 : _GEN_1637; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1639 = 8'h67 == _t_T_10[31:24] ? 8'h85 : _GEN_1638; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1640 = 8'h68 == _t_T_10[31:24] ? 8'h45 : _GEN_1639; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1641 = 8'h69 == _t_T_10[31:24] ? 8'hf9 : _GEN_1640; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1642 = 8'h6a == _t_T_10[31:24] ? 8'h2 : _GEN_1641; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1643 = 8'h6b == _t_T_10[31:24] ? 8'h7f : _GEN_1642; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1644 = 8'h6c == _t_T_10[31:24] ? 8'h50 : _GEN_1643; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1645 = 8'h6d == _t_T_10[31:24] ? 8'h3c : _GEN_1644; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1646 = 8'h6e == _t_T_10[31:24] ? 8'h9f : _GEN_1645; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1647 = 8'h6f == _t_T_10[31:24] ? 8'ha8 : _GEN_1646; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1648 = 8'h70 == _t_T_10[31:24] ? 8'h51 : _GEN_1647; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1649 = 8'h71 == _t_T_10[31:24] ? 8'ha3 : _GEN_1648; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1650 = 8'h72 == _t_T_10[31:24] ? 8'h40 : _GEN_1649; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1651 = 8'h73 == _t_T_10[31:24] ? 8'h8f : _GEN_1650; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1652 = 8'h74 == _t_T_10[31:24] ? 8'h92 : _GEN_1651; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1653 = 8'h75 == _t_T_10[31:24] ? 8'h9d : _GEN_1652; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1654 = 8'h76 == _t_T_10[31:24] ? 8'h38 : _GEN_1653; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1655 = 8'h77 == _t_T_10[31:24] ? 8'hf5 : _GEN_1654; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1656 = 8'h78 == _t_T_10[31:24] ? 8'hbc : _GEN_1655; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1657 = 8'h79 == _t_T_10[31:24] ? 8'hb6 : _GEN_1656; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1658 = 8'h7a == _t_T_10[31:24] ? 8'hda : _GEN_1657; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1659 = 8'h7b == _t_T_10[31:24] ? 8'h21 : _GEN_1658; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1660 = 8'h7c == _t_T_10[31:24] ? 8'h10 : _GEN_1659; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1661 = 8'h7d == _t_T_10[31:24] ? 8'hff : _GEN_1660; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1662 = 8'h7e == _t_T_10[31:24] ? 8'hf3 : _GEN_1661; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1663 = 8'h7f == _t_T_10[31:24] ? 8'hd2 : _GEN_1662; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1664 = 8'h80 == _t_T_10[31:24] ? 8'hcd : _GEN_1663; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1665 = 8'h81 == _t_T_10[31:24] ? 8'hc : _GEN_1664; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1666 = 8'h82 == _t_T_10[31:24] ? 8'h13 : _GEN_1665; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1667 = 8'h83 == _t_T_10[31:24] ? 8'hec : _GEN_1666; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1668 = 8'h84 == _t_T_10[31:24] ? 8'h5f : _GEN_1667; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1669 = 8'h85 == _t_T_10[31:24] ? 8'h97 : _GEN_1668; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1670 = 8'h86 == _t_T_10[31:24] ? 8'h44 : _GEN_1669; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1671 = 8'h87 == _t_T_10[31:24] ? 8'h17 : _GEN_1670; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1672 = 8'h88 == _t_T_10[31:24] ? 8'hc4 : _GEN_1671; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1673 = 8'h89 == _t_T_10[31:24] ? 8'ha7 : _GEN_1672; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1674 = 8'h8a == _t_T_10[31:24] ? 8'h7e : _GEN_1673; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1675 = 8'h8b == _t_T_10[31:24] ? 8'h3d : _GEN_1674; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1676 = 8'h8c == _t_T_10[31:24] ? 8'h64 : _GEN_1675; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1677 = 8'h8d == _t_T_10[31:24] ? 8'h5d : _GEN_1676; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1678 = 8'h8e == _t_T_10[31:24] ? 8'h19 : _GEN_1677; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1679 = 8'h8f == _t_T_10[31:24] ? 8'h73 : _GEN_1678; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1680 = 8'h90 == _t_T_10[31:24] ? 8'h60 : _GEN_1679; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1681 = 8'h91 == _t_T_10[31:24] ? 8'h81 : _GEN_1680; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1682 = 8'h92 == _t_T_10[31:24] ? 8'h4f : _GEN_1681; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1683 = 8'h93 == _t_T_10[31:24] ? 8'hdc : _GEN_1682; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1684 = 8'h94 == _t_T_10[31:24] ? 8'h22 : _GEN_1683; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1685 = 8'h95 == _t_T_10[31:24] ? 8'h2a : _GEN_1684; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1686 = 8'h96 == _t_T_10[31:24] ? 8'h90 : _GEN_1685; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1687 = 8'h97 == _t_T_10[31:24] ? 8'h88 : _GEN_1686; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1688 = 8'h98 == _t_T_10[31:24] ? 8'h46 : _GEN_1687; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1689 = 8'h99 == _t_T_10[31:24] ? 8'hee : _GEN_1688; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1690 = 8'h9a == _t_T_10[31:24] ? 8'hb8 : _GEN_1689; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1691 = 8'h9b == _t_T_10[31:24] ? 8'h14 : _GEN_1690; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1692 = 8'h9c == _t_T_10[31:24] ? 8'hde : _GEN_1691; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1693 = 8'h9d == _t_T_10[31:24] ? 8'h5e : _GEN_1692; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1694 = 8'h9e == _t_T_10[31:24] ? 8'hb : _GEN_1693; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1695 = 8'h9f == _t_T_10[31:24] ? 8'hdb : _GEN_1694; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1696 = 8'ha0 == _t_T_10[31:24] ? 8'he0 : _GEN_1695; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1697 = 8'ha1 == _t_T_10[31:24] ? 8'h32 : _GEN_1696; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1698 = 8'ha2 == _t_T_10[31:24] ? 8'h3a : _GEN_1697; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1699 = 8'ha3 == _t_T_10[31:24] ? 8'ha : _GEN_1698; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1700 = 8'ha4 == _t_T_10[31:24] ? 8'h49 : _GEN_1699; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1701 = 8'ha5 == _t_T_10[31:24] ? 8'h6 : _GEN_1700; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1702 = 8'ha6 == _t_T_10[31:24] ? 8'h24 : _GEN_1701; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1703 = 8'ha7 == _t_T_10[31:24] ? 8'h5c : _GEN_1702; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1704 = 8'ha8 == _t_T_10[31:24] ? 8'hc2 : _GEN_1703; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1705 = 8'ha9 == _t_T_10[31:24] ? 8'hd3 : _GEN_1704; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1706 = 8'haa == _t_T_10[31:24] ? 8'hac : _GEN_1705; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1707 = 8'hab == _t_T_10[31:24] ? 8'h62 : _GEN_1706; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1708 = 8'hac == _t_T_10[31:24] ? 8'h91 : _GEN_1707; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1709 = 8'had == _t_T_10[31:24] ? 8'h95 : _GEN_1708; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1710 = 8'hae == _t_T_10[31:24] ? 8'he4 : _GEN_1709; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1711 = 8'haf == _t_T_10[31:24] ? 8'h79 : _GEN_1710; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1712 = 8'hb0 == _t_T_10[31:24] ? 8'he7 : _GEN_1711; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1713 = 8'hb1 == _t_T_10[31:24] ? 8'hc8 : _GEN_1712; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1714 = 8'hb2 == _t_T_10[31:24] ? 8'h37 : _GEN_1713; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1715 = 8'hb3 == _t_T_10[31:24] ? 8'h6d : _GEN_1714; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1716 = 8'hb4 == _t_T_10[31:24] ? 8'h8d : _GEN_1715; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1717 = 8'hb5 == _t_T_10[31:24] ? 8'hd5 : _GEN_1716; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1718 = 8'hb6 == _t_T_10[31:24] ? 8'h4e : _GEN_1717; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1719 = 8'hb7 == _t_T_10[31:24] ? 8'ha9 : _GEN_1718; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1720 = 8'hb8 == _t_T_10[31:24] ? 8'h6c : _GEN_1719; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1721 = 8'hb9 == _t_T_10[31:24] ? 8'h56 : _GEN_1720; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1722 = 8'hba == _t_T_10[31:24] ? 8'hf4 : _GEN_1721; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1723 = 8'hbb == _t_T_10[31:24] ? 8'hea : _GEN_1722; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1724 = 8'hbc == _t_T_10[31:24] ? 8'h65 : _GEN_1723; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1725 = 8'hbd == _t_T_10[31:24] ? 8'h7a : _GEN_1724; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1726 = 8'hbe == _t_T_10[31:24] ? 8'hae : _GEN_1725; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1727 = 8'hbf == _t_T_10[31:24] ? 8'h8 : _GEN_1726; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1728 = 8'hc0 == _t_T_10[31:24] ? 8'hba : _GEN_1727; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1729 = 8'hc1 == _t_T_10[31:24] ? 8'h78 : _GEN_1728; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1730 = 8'hc2 == _t_T_10[31:24] ? 8'h25 : _GEN_1729; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1731 = 8'hc3 == _t_T_10[31:24] ? 8'h2e : _GEN_1730; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1732 = 8'hc4 == _t_T_10[31:24] ? 8'h1c : _GEN_1731; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1733 = 8'hc5 == _t_T_10[31:24] ? 8'ha6 : _GEN_1732; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1734 = 8'hc6 == _t_T_10[31:24] ? 8'hb4 : _GEN_1733; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1735 = 8'hc7 == _t_T_10[31:24] ? 8'hc6 : _GEN_1734; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1736 = 8'hc8 == _t_T_10[31:24] ? 8'he8 : _GEN_1735; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1737 = 8'hc9 == _t_T_10[31:24] ? 8'hdd : _GEN_1736; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1738 = 8'hca == _t_T_10[31:24] ? 8'h74 : _GEN_1737; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1739 = 8'hcb == _t_T_10[31:24] ? 8'h1f : _GEN_1738; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1740 = 8'hcc == _t_T_10[31:24] ? 8'h4b : _GEN_1739; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1741 = 8'hcd == _t_T_10[31:24] ? 8'hbd : _GEN_1740; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1742 = 8'hce == _t_T_10[31:24] ? 8'h8b : _GEN_1741; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1743 = 8'hcf == _t_T_10[31:24] ? 8'h8a : _GEN_1742; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1744 = 8'hd0 == _t_T_10[31:24] ? 8'h70 : _GEN_1743; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1745 = 8'hd1 == _t_T_10[31:24] ? 8'h3e : _GEN_1744; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1746 = 8'hd2 == _t_T_10[31:24] ? 8'hb5 : _GEN_1745; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1747 = 8'hd3 == _t_T_10[31:24] ? 8'h66 : _GEN_1746; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1748 = 8'hd4 == _t_T_10[31:24] ? 8'h48 : _GEN_1747; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1749 = 8'hd5 == _t_T_10[31:24] ? 8'h3 : _GEN_1748; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1750 = 8'hd6 == _t_T_10[31:24] ? 8'hf6 : _GEN_1749; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1751 = 8'hd7 == _t_T_10[31:24] ? 8'he : _GEN_1750; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1752 = 8'hd8 == _t_T_10[31:24] ? 8'h61 : _GEN_1751; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1753 = 8'hd9 == _t_T_10[31:24] ? 8'h35 : _GEN_1752; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1754 = 8'hda == _t_T_10[31:24] ? 8'h57 : _GEN_1753; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1755 = 8'hdb == _t_T_10[31:24] ? 8'hb9 : _GEN_1754; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1756 = 8'hdc == _t_T_10[31:24] ? 8'h86 : _GEN_1755; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1757 = 8'hdd == _t_T_10[31:24] ? 8'hc1 : _GEN_1756; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1758 = 8'hde == _t_T_10[31:24] ? 8'h1d : _GEN_1757; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1759 = 8'hdf == _t_T_10[31:24] ? 8'h9e : _GEN_1758; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1760 = 8'he0 == _t_T_10[31:24] ? 8'he1 : _GEN_1759; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1761 = 8'he1 == _t_T_10[31:24] ? 8'hf8 : _GEN_1760; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1762 = 8'he2 == _t_T_10[31:24] ? 8'h98 : _GEN_1761; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1763 = 8'he3 == _t_T_10[31:24] ? 8'h11 : _GEN_1762; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1764 = 8'he4 == _t_T_10[31:24] ? 8'h69 : _GEN_1763; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1765 = 8'he5 == _t_T_10[31:24] ? 8'hd9 : _GEN_1764; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1766 = 8'he6 == _t_T_10[31:24] ? 8'h8e : _GEN_1765; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1767 = 8'he7 == _t_T_10[31:24] ? 8'h94 : _GEN_1766; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1768 = 8'he8 == _t_T_10[31:24] ? 8'h9b : _GEN_1767; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1769 = 8'he9 == _t_T_10[31:24] ? 8'h1e : _GEN_1768; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1770 = 8'hea == _t_T_10[31:24] ? 8'h87 : _GEN_1769; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1771 = 8'heb == _t_T_10[31:24] ? 8'he9 : _GEN_1770; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1772 = 8'hec == _t_T_10[31:24] ? 8'hce : _GEN_1771; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1773 = 8'hed == _t_T_10[31:24] ? 8'h55 : _GEN_1772; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1774 = 8'hee == _t_T_10[31:24] ? 8'h28 : _GEN_1773; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1775 = 8'hef == _t_T_10[31:24] ? 8'hdf : _GEN_1774; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1776 = 8'hf0 == _t_T_10[31:24] ? 8'h8c : _GEN_1775; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1777 = 8'hf1 == _t_T_10[31:24] ? 8'ha1 : _GEN_1776; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1778 = 8'hf2 == _t_T_10[31:24] ? 8'h89 : _GEN_1777; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1779 = 8'hf3 == _t_T_10[31:24] ? 8'hd : _GEN_1778; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1780 = 8'hf4 == _t_T_10[31:24] ? 8'hbf : _GEN_1779; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1781 = 8'hf5 == _t_T_10[31:24] ? 8'he6 : _GEN_1780; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1782 = 8'hf6 == _t_T_10[31:24] ? 8'h42 : _GEN_1781; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1783 = 8'hf7 == _t_T_10[31:24] ? 8'h68 : _GEN_1782; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1784 = 8'hf8 == _t_T_10[31:24] ? 8'h41 : _GEN_1783; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1785 = 8'hf9 == _t_T_10[31:24] ? 8'h99 : _GEN_1784; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1786 = 8'hfa == _t_T_10[31:24] ? 8'h2d : _GEN_1785; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1787 = 8'hfb == _t_T_10[31:24] ? 8'hf : _GEN_1786; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1788 = 8'hfc == _t_T_10[31:24] ? 8'hb0 : _GEN_1787; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1789 = 8'hfd == _t_T_10[31:24] ? 8'h54 : _GEN_1788; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1790 = 8'hfe == _t_T_10[31:24] ? 8'hbb : _GEN_1789; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1791 = 8'hff == _t_T_10[31:24] ? 8'h16 : _GEN_1790; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1793 = 8'h1 == _t_T_10[23:16] ? 8'h7c : 8'h63; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1794 = 8'h2 == _t_T_10[23:16] ? 8'h77 : _GEN_1793; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1795 = 8'h3 == _t_T_10[23:16] ? 8'h7b : _GEN_1794; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1796 = 8'h4 == _t_T_10[23:16] ? 8'hf2 : _GEN_1795; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1797 = 8'h5 == _t_T_10[23:16] ? 8'h6b : _GEN_1796; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1798 = 8'h6 == _t_T_10[23:16] ? 8'h6f : _GEN_1797; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1799 = 8'h7 == _t_T_10[23:16] ? 8'hc5 : _GEN_1798; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1800 = 8'h8 == _t_T_10[23:16] ? 8'h30 : _GEN_1799; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1801 = 8'h9 == _t_T_10[23:16] ? 8'h1 : _GEN_1800; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1802 = 8'ha == _t_T_10[23:16] ? 8'h67 : _GEN_1801; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1803 = 8'hb == _t_T_10[23:16] ? 8'h2b : _GEN_1802; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1804 = 8'hc == _t_T_10[23:16] ? 8'hfe : _GEN_1803; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1805 = 8'hd == _t_T_10[23:16] ? 8'hd7 : _GEN_1804; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1806 = 8'he == _t_T_10[23:16] ? 8'hab : _GEN_1805; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1807 = 8'hf == _t_T_10[23:16] ? 8'h76 : _GEN_1806; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1808 = 8'h10 == _t_T_10[23:16] ? 8'hca : _GEN_1807; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1809 = 8'h11 == _t_T_10[23:16] ? 8'h82 : _GEN_1808; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1810 = 8'h12 == _t_T_10[23:16] ? 8'hc9 : _GEN_1809; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1811 = 8'h13 == _t_T_10[23:16] ? 8'h7d : _GEN_1810; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1812 = 8'h14 == _t_T_10[23:16] ? 8'hfa : _GEN_1811; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1813 = 8'h15 == _t_T_10[23:16] ? 8'h59 : _GEN_1812; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1814 = 8'h16 == _t_T_10[23:16] ? 8'h47 : _GEN_1813; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1815 = 8'h17 == _t_T_10[23:16] ? 8'hf0 : _GEN_1814; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1816 = 8'h18 == _t_T_10[23:16] ? 8'had : _GEN_1815; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1817 = 8'h19 == _t_T_10[23:16] ? 8'hd4 : _GEN_1816; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1818 = 8'h1a == _t_T_10[23:16] ? 8'ha2 : _GEN_1817; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1819 = 8'h1b == _t_T_10[23:16] ? 8'haf : _GEN_1818; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1820 = 8'h1c == _t_T_10[23:16] ? 8'h9c : _GEN_1819; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1821 = 8'h1d == _t_T_10[23:16] ? 8'ha4 : _GEN_1820; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1822 = 8'h1e == _t_T_10[23:16] ? 8'h72 : _GEN_1821; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1823 = 8'h1f == _t_T_10[23:16] ? 8'hc0 : _GEN_1822; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1824 = 8'h20 == _t_T_10[23:16] ? 8'hb7 : _GEN_1823; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1825 = 8'h21 == _t_T_10[23:16] ? 8'hfd : _GEN_1824; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1826 = 8'h22 == _t_T_10[23:16] ? 8'h93 : _GEN_1825; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1827 = 8'h23 == _t_T_10[23:16] ? 8'h26 : _GEN_1826; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1828 = 8'h24 == _t_T_10[23:16] ? 8'h36 : _GEN_1827; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1829 = 8'h25 == _t_T_10[23:16] ? 8'h3f : _GEN_1828; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1830 = 8'h26 == _t_T_10[23:16] ? 8'hf7 : _GEN_1829; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1831 = 8'h27 == _t_T_10[23:16] ? 8'hcc : _GEN_1830; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1832 = 8'h28 == _t_T_10[23:16] ? 8'h34 : _GEN_1831; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1833 = 8'h29 == _t_T_10[23:16] ? 8'ha5 : _GEN_1832; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1834 = 8'h2a == _t_T_10[23:16] ? 8'he5 : _GEN_1833; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1835 = 8'h2b == _t_T_10[23:16] ? 8'hf1 : _GEN_1834; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1836 = 8'h2c == _t_T_10[23:16] ? 8'h71 : _GEN_1835; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1837 = 8'h2d == _t_T_10[23:16] ? 8'hd8 : _GEN_1836; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1838 = 8'h2e == _t_T_10[23:16] ? 8'h31 : _GEN_1837; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1839 = 8'h2f == _t_T_10[23:16] ? 8'h15 : _GEN_1838; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1840 = 8'h30 == _t_T_10[23:16] ? 8'h4 : _GEN_1839; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1841 = 8'h31 == _t_T_10[23:16] ? 8'hc7 : _GEN_1840; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1842 = 8'h32 == _t_T_10[23:16] ? 8'h23 : _GEN_1841; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1843 = 8'h33 == _t_T_10[23:16] ? 8'hc3 : _GEN_1842; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1844 = 8'h34 == _t_T_10[23:16] ? 8'h18 : _GEN_1843; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1845 = 8'h35 == _t_T_10[23:16] ? 8'h96 : _GEN_1844; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1846 = 8'h36 == _t_T_10[23:16] ? 8'h5 : _GEN_1845; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1847 = 8'h37 == _t_T_10[23:16] ? 8'h9a : _GEN_1846; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1848 = 8'h38 == _t_T_10[23:16] ? 8'h7 : _GEN_1847; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1849 = 8'h39 == _t_T_10[23:16] ? 8'h12 : _GEN_1848; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1850 = 8'h3a == _t_T_10[23:16] ? 8'h80 : _GEN_1849; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1851 = 8'h3b == _t_T_10[23:16] ? 8'he2 : _GEN_1850; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1852 = 8'h3c == _t_T_10[23:16] ? 8'heb : _GEN_1851; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1853 = 8'h3d == _t_T_10[23:16] ? 8'h27 : _GEN_1852; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1854 = 8'h3e == _t_T_10[23:16] ? 8'hb2 : _GEN_1853; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1855 = 8'h3f == _t_T_10[23:16] ? 8'h75 : _GEN_1854; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1856 = 8'h40 == _t_T_10[23:16] ? 8'h9 : _GEN_1855; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1857 = 8'h41 == _t_T_10[23:16] ? 8'h83 : _GEN_1856; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1858 = 8'h42 == _t_T_10[23:16] ? 8'h2c : _GEN_1857; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1859 = 8'h43 == _t_T_10[23:16] ? 8'h1a : _GEN_1858; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1860 = 8'h44 == _t_T_10[23:16] ? 8'h1b : _GEN_1859; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1861 = 8'h45 == _t_T_10[23:16] ? 8'h6e : _GEN_1860; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1862 = 8'h46 == _t_T_10[23:16] ? 8'h5a : _GEN_1861; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1863 = 8'h47 == _t_T_10[23:16] ? 8'ha0 : _GEN_1862; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1864 = 8'h48 == _t_T_10[23:16] ? 8'h52 : _GEN_1863; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1865 = 8'h49 == _t_T_10[23:16] ? 8'h3b : _GEN_1864; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1866 = 8'h4a == _t_T_10[23:16] ? 8'hd6 : _GEN_1865; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1867 = 8'h4b == _t_T_10[23:16] ? 8'hb3 : _GEN_1866; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1868 = 8'h4c == _t_T_10[23:16] ? 8'h29 : _GEN_1867; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1869 = 8'h4d == _t_T_10[23:16] ? 8'he3 : _GEN_1868; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1870 = 8'h4e == _t_T_10[23:16] ? 8'h2f : _GEN_1869; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1871 = 8'h4f == _t_T_10[23:16] ? 8'h84 : _GEN_1870; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1872 = 8'h50 == _t_T_10[23:16] ? 8'h53 : _GEN_1871; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1873 = 8'h51 == _t_T_10[23:16] ? 8'hd1 : _GEN_1872; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1874 = 8'h52 == _t_T_10[23:16] ? 8'h0 : _GEN_1873; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1875 = 8'h53 == _t_T_10[23:16] ? 8'hed : _GEN_1874; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1876 = 8'h54 == _t_T_10[23:16] ? 8'h20 : _GEN_1875; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1877 = 8'h55 == _t_T_10[23:16] ? 8'hfc : _GEN_1876; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1878 = 8'h56 == _t_T_10[23:16] ? 8'hb1 : _GEN_1877; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1879 = 8'h57 == _t_T_10[23:16] ? 8'h5b : _GEN_1878; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1880 = 8'h58 == _t_T_10[23:16] ? 8'h6a : _GEN_1879; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1881 = 8'h59 == _t_T_10[23:16] ? 8'hcb : _GEN_1880; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1882 = 8'h5a == _t_T_10[23:16] ? 8'hbe : _GEN_1881; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1883 = 8'h5b == _t_T_10[23:16] ? 8'h39 : _GEN_1882; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1884 = 8'h5c == _t_T_10[23:16] ? 8'h4a : _GEN_1883; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1885 = 8'h5d == _t_T_10[23:16] ? 8'h4c : _GEN_1884; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1886 = 8'h5e == _t_T_10[23:16] ? 8'h58 : _GEN_1885; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1887 = 8'h5f == _t_T_10[23:16] ? 8'hcf : _GEN_1886; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1888 = 8'h60 == _t_T_10[23:16] ? 8'hd0 : _GEN_1887; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1889 = 8'h61 == _t_T_10[23:16] ? 8'hef : _GEN_1888; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1890 = 8'h62 == _t_T_10[23:16] ? 8'haa : _GEN_1889; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1891 = 8'h63 == _t_T_10[23:16] ? 8'hfb : _GEN_1890; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1892 = 8'h64 == _t_T_10[23:16] ? 8'h43 : _GEN_1891; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1893 = 8'h65 == _t_T_10[23:16] ? 8'h4d : _GEN_1892; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1894 = 8'h66 == _t_T_10[23:16] ? 8'h33 : _GEN_1893; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1895 = 8'h67 == _t_T_10[23:16] ? 8'h85 : _GEN_1894; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1896 = 8'h68 == _t_T_10[23:16] ? 8'h45 : _GEN_1895; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1897 = 8'h69 == _t_T_10[23:16] ? 8'hf9 : _GEN_1896; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1898 = 8'h6a == _t_T_10[23:16] ? 8'h2 : _GEN_1897; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1899 = 8'h6b == _t_T_10[23:16] ? 8'h7f : _GEN_1898; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1900 = 8'h6c == _t_T_10[23:16] ? 8'h50 : _GEN_1899; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1901 = 8'h6d == _t_T_10[23:16] ? 8'h3c : _GEN_1900; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1902 = 8'h6e == _t_T_10[23:16] ? 8'h9f : _GEN_1901; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1903 = 8'h6f == _t_T_10[23:16] ? 8'ha8 : _GEN_1902; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1904 = 8'h70 == _t_T_10[23:16] ? 8'h51 : _GEN_1903; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1905 = 8'h71 == _t_T_10[23:16] ? 8'ha3 : _GEN_1904; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1906 = 8'h72 == _t_T_10[23:16] ? 8'h40 : _GEN_1905; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1907 = 8'h73 == _t_T_10[23:16] ? 8'h8f : _GEN_1906; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1908 = 8'h74 == _t_T_10[23:16] ? 8'h92 : _GEN_1907; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1909 = 8'h75 == _t_T_10[23:16] ? 8'h9d : _GEN_1908; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1910 = 8'h76 == _t_T_10[23:16] ? 8'h38 : _GEN_1909; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1911 = 8'h77 == _t_T_10[23:16] ? 8'hf5 : _GEN_1910; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1912 = 8'h78 == _t_T_10[23:16] ? 8'hbc : _GEN_1911; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1913 = 8'h79 == _t_T_10[23:16] ? 8'hb6 : _GEN_1912; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1914 = 8'h7a == _t_T_10[23:16] ? 8'hda : _GEN_1913; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1915 = 8'h7b == _t_T_10[23:16] ? 8'h21 : _GEN_1914; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1916 = 8'h7c == _t_T_10[23:16] ? 8'h10 : _GEN_1915; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1917 = 8'h7d == _t_T_10[23:16] ? 8'hff : _GEN_1916; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1918 = 8'h7e == _t_T_10[23:16] ? 8'hf3 : _GEN_1917; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1919 = 8'h7f == _t_T_10[23:16] ? 8'hd2 : _GEN_1918; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1920 = 8'h80 == _t_T_10[23:16] ? 8'hcd : _GEN_1919; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1921 = 8'h81 == _t_T_10[23:16] ? 8'hc : _GEN_1920; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1922 = 8'h82 == _t_T_10[23:16] ? 8'h13 : _GEN_1921; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1923 = 8'h83 == _t_T_10[23:16] ? 8'hec : _GEN_1922; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1924 = 8'h84 == _t_T_10[23:16] ? 8'h5f : _GEN_1923; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1925 = 8'h85 == _t_T_10[23:16] ? 8'h97 : _GEN_1924; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1926 = 8'h86 == _t_T_10[23:16] ? 8'h44 : _GEN_1925; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1927 = 8'h87 == _t_T_10[23:16] ? 8'h17 : _GEN_1926; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1928 = 8'h88 == _t_T_10[23:16] ? 8'hc4 : _GEN_1927; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1929 = 8'h89 == _t_T_10[23:16] ? 8'ha7 : _GEN_1928; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1930 = 8'h8a == _t_T_10[23:16] ? 8'h7e : _GEN_1929; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1931 = 8'h8b == _t_T_10[23:16] ? 8'h3d : _GEN_1930; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1932 = 8'h8c == _t_T_10[23:16] ? 8'h64 : _GEN_1931; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1933 = 8'h8d == _t_T_10[23:16] ? 8'h5d : _GEN_1932; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1934 = 8'h8e == _t_T_10[23:16] ? 8'h19 : _GEN_1933; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1935 = 8'h8f == _t_T_10[23:16] ? 8'h73 : _GEN_1934; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1936 = 8'h90 == _t_T_10[23:16] ? 8'h60 : _GEN_1935; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1937 = 8'h91 == _t_T_10[23:16] ? 8'h81 : _GEN_1936; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1938 = 8'h92 == _t_T_10[23:16] ? 8'h4f : _GEN_1937; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1939 = 8'h93 == _t_T_10[23:16] ? 8'hdc : _GEN_1938; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1940 = 8'h94 == _t_T_10[23:16] ? 8'h22 : _GEN_1939; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1941 = 8'h95 == _t_T_10[23:16] ? 8'h2a : _GEN_1940; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1942 = 8'h96 == _t_T_10[23:16] ? 8'h90 : _GEN_1941; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1943 = 8'h97 == _t_T_10[23:16] ? 8'h88 : _GEN_1942; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1944 = 8'h98 == _t_T_10[23:16] ? 8'h46 : _GEN_1943; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1945 = 8'h99 == _t_T_10[23:16] ? 8'hee : _GEN_1944; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1946 = 8'h9a == _t_T_10[23:16] ? 8'hb8 : _GEN_1945; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1947 = 8'h9b == _t_T_10[23:16] ? 8'h14 : _GEN_1946; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1948 = 8'h9c == _t_T_10[23:16] ? 8'hde : _GEN_1947; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1949 = 8'h9d == _t_T_10[23:16] ? 8'h5e : _GEN_1948; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1950 = 8'h9e == _t_T_10[23:16] ? 8'hb : _GEN_1949; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1951 = 8'h9f == _t_T_10[23:16] ? 8'hdb : _GEN_1950; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1952 = 8'ha0 == _t_T_10[23:16] ? 8'he0 : _GEN_1951; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1953 = 8'ha1 == _t_T_10[23:16] ? 8'h32 : _GEN_1952; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1954 = 8'ha2 == _t_T_10[23:16] ? 8'h3a : _GEN_1953; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1955 = 8'ha3 == _t_T_10[23:16] ? 8'ha : _GEN_1954; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1956 = 8'ha4 == _t_T_10[23:16] ? 8'h49 : _GEN_1955; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1957 = 8'ha5 == _t_T_10[23:16] ? 8'h6 : _GEN_1956; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1958 = 8'ha6 == _t_T_10[23:16] ? 8'h24 : _GEN_1957; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1959 = 8'ha7 == _t_T_10[23:16] ? 8'h5c : _GEN_1958; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1960 = 8'ha8 == _t_T_10[23:16] ? 8'hc2 : _GEN_1959; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1961 = 8'ha9 == _t_T_10[23:16] ? 8'hd3 : _GEN_1960; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1962 = 8'haa == _t_T_10[23:16] ? 8'hac : _GEN_1961; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1963 = 8'hab == _t_T_10[23:16] ? 8'h62 : _GEN_1962; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1964 = 8'hac == _t_T_10[23:16] ? 8'h91 : _GEN_1963; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1965 = 8'had == _t_T_10[23:16] ? 8'h95 : _GEN_1964; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1966 = 8'hae == _t_T_10[23:16] ? 8'he4 : _GEN_1965; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1967 = 8'haf == _t_T_10[23:16] ? 8'h79 : _GEN_1966; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1968 = 8'hb0 == _t_T_10[23:16] ? 8'he7 : _GEN_1967; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1969 = 8'hb1 == _t_T_10[23:16] ? 8'hc8 : _GEN_1968; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1970 = 8'hb2 == _t_T_10[23:16] ? 8'h37 : _GEN_1969; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1971 = 8'hb3 == _t_T_10[23:16] ? 8'h6d : _GEN_1970; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1972 = 8'hb4 == _t_T_10[23:16] ? 8'h8d : _GEN_1971; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1973 = 8'hb5 == _t_T_10[23:16] ? 8'hd5 : _GEN_1972; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1974 = 8'hb6 == _t_T_10[23:16] ? 8'h4e : _GEN_1973; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1975 = 8'hb7 == _t_T_10[23:16] ? 8'ha9 : _GEN_1974; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1976 = 8'hb8 == _t_T_10[23:16] ? 8'h6c : _GEN_1975; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1977 = 8'hb9 == _t_T_10[23:16] ? 8'h56 : _GEN_1976; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1978 = 8'hba == _t_T_10[23:16] ? 8'hf4 : _GEN_1977; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1979 = 8'hbb == _t_T_10[23:16] ? 8'hea : _GEN_1978; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1980 = 8'hbc == _t_T_10[23:16] ? 8'h65 : _GEN_1979; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1981 = 8'hbd == _t_T_10[23:16] ? 8'h7a : _GEN_1980; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1982 = 8'hbe == _t_T_10[23:16] ? 8'hae : _GEN_1981; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1983 = 8'hbf == _t_T_10[23:16] ? 8'h8 : _GEN_1982; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1984 = 8'hc0 == _t_T_10[23:16] ? 8'hba : _GEN_1983; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1985 = 8'hc1 == _t_T_10[23:16] ? 8'h78 : _GEN_1984; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1986 = 8'hc2 == _t_T_10[23:16] ? 8'h25 : _GEN_1985; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1987 = 8'hc3 == _t_T_10[23:16] ? 8'h2e : _GEN_1986; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1988 = 8'hc4 == _t_T_10[23:16] ? 8'h1c : _GEN_1987; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1989 = 8'hc5 == _t_T_10[23:16] ? 8'ha6 : _GEN_1988; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1990 = 8'hc6 == _t_T_10[23:16] ? 8'hb4 : _GEN_1989; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1991 = 8'hc7 == _t_T_10[23:16] ? 8'hc6 : _GEN_1990; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1992 = 8'hc8 == _t_T_10[23:16] ? 8'he8 : _GEN_1991; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1993 = 8'hc9 == _t_T_10[23:16] ? 8'hdd : _GEN_1992; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1994 = 8'hca == _t_T_10[23:16] ? 8'h74 : _GEN_1993; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1995 = 8'hcb == _t_T_10[23:16] ? 8'h1f : _GEN_1994; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1996 = 8'hcc == _t_T_10[23:16] ? 8'h4b : _GEN_1995; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1997 = 8'hcd == _t_T_10[23:16] ? 8'hbd : _GEN_1996; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1998 = 8'hce == _t_T_10[23:16] ? 8'h8b : _GEN_1997; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_1999 = 8'hcf == _t_T_10[23:16] ? 8'h8a : _GEN_1998; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2000 = 8'hd0 == _t_T_10[23:16] ? 8'h70 : _GEN_1999; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2001 = 8'hd1 == _t_T_10[23:16] ? 8'h3e : _GEN_2000; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2002 = 8'hd2 == _t_T_10[23:16] ? 8'hb5 : _GEN_2001; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2003 = 8'hd3 == _t_T_10[23:16] ? 8'h66 : _GEN_2002; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2004 = 8'hd4 == _t_T_10[23:16] ? 8'h48 : _GEN_2003; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2005 = 8'hd5 == _t_T_10[23:16] ? 8'h3 : _GEN_2004; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2006 = 8'hd6 == _t_T_10[23:16] ? 8'hf6 : _GEN_2005; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2007 = 8'hd7 == _t_T_10[23:16] ? 8'he : _GEN_2006; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2008 = 8'hd8 == _t_T_10[23:16] ? 8'h61 : _GEN_2007; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2009 = 8'hd9 == _t_T_10[23:16] ? 8'h35 : _GEN_2008; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2010 = 8'hda == _t_T_10[23:16] ? 8'h57 : _GEN_2009; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2011 = 8'hdb == _t_T_10[23:16] ? 8'hb9 : _GEN_2010; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2012 = 8'hdc == _t_T_10[23:16] ? 8'h86 : _GEN_2011; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2013 = 8'hdd == _t_T_10[23:16] ? 8'hc1 : _GEN_2012; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2014 = 8'hde == _t_T_10[23:16] ? 8'h1d : _GEN_2013; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2015 = 8'hdf == _t_T_10[23:16] ? 8'h9e : _GEN_2014; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2016 = 8'he0 == _t_T_10[23:16] ? 8'he1 : _GEN_2015; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2017 = 8'he1 == _t_T_10[23:16] ? 8'hf8 : _GEN_2016; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2018 = 8'he2 == _t_T_10[23:16] ? 8'h98 : _GEN_2017; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2019 = 8'he3 == _t_T_10[23:16] ? 8'h11 : _GEN_2018; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2020 = 8'he4 == _t_T_10[23:16] ? 8'h69 : _GEN_2019; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2021 = 8'he5 == _t_T_10[23:16] ? 8'hd9 : _GEN_2020; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2022 = 8'he6 == _t_T_10[23:16] ? 8'h8e : _GEN_2021; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2023 = 8'he7 == _t_T_10[23:16] ? 8'h94 : _GEN_2022; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2024 = 8'he8 == _t_T_10[23:16] ? 8'h9b : _GEN_2023; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2025 = 8'he9 == _t_T_10[23:16] ? 8'h1e : _GEN_2024; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2026 = 8'hea == _t_T_10[23:16] ? 8'h87 : _GEN_2025; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2027 = 8'heb == _t_T_10[23:16] ? 8'he9 : _GEN_2026; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2028 = 8'hec == _t_T_10[23:16] ? 8'hce : _GEN_2027; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2029 = 8'hed == _t_T_10[23:16] ? 8'h55 : _GEN_2028; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2030 = 8'hee == _t_T_10[23:16] ? 8'h28 : _GEN_2029; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2031 = 8'hef == _t_T_10[23:16] ? 8'hdf : _GEN_2030; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2032 = 8'hf0 == _t_T_10[23:16] ? 8'h8c : _GEN_2031; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2033 = 8'hf1 == _t_T_10[23:16] ? 8'ha1 : _GEN_2032; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2034 = 8'hf2 == _t_T_10[23:16] ? 8'h89 : _GEN_2033; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2035 = 8'hf3 == _t_T_10[23:16] ? 8'hd : _GEN_2034; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2036 = 8'hf4 == _t_T_10[23:16] ? 8'hbf : _GEN_2035; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2037 = 8'hf5 == _t_T_10[23:16] ? 8'he6 : _GEN_2036; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2038 = 8'hf6 == _t_T_10[23:16] ? 8'h42 : _GEN_2037; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2039 = 8'hf7 == _t_T_10[23:16] ? 8'h68 : _GEN_2038; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2040 = 8'hf8 == _t_T_10[23:16] ? 8'h41 : _GEN_2039; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2041 = 8'hf9 == _t_T_10[23:16] ? 8'h99 : _GEN_2040; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2042 = 8'hfa == _t_T_10[23:16] ? 8'h2d : _GEN_2041; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2043 = 8'hfb == _t_T_10[23:16] ? 8'hf : _GEN_2042; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2044 = 8'hfc == _t_T_10[23:16] ? 8'hb0 : _GEN_2043; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2045 = 8'hfd == _t_T_10[23:16] ? 8'h54 : _GEN_2044; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2046 = 8'hfe == _t_T_10[23:16] ? 8'hbb : _GEN_2045; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2047 = 8'hff == _t_T_10[23:16] ? 8'h16 : _GEN_2046; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [31:0] _t_T_15 = {_GEN_1791,_GEN_2047,_GEN_1279,_GEN_1535}; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:8]
  wire [31:0] t_1 = _t_T_15 ^ 32'h2000000; // @[src/main/scala/crypto/aes/KeySchedule.scala 59:32]
  wire [31:0] w_8 = w_4 ^ t_1; // @[src/main/scala/crypto/aes/KeySchedule.scala 63:21]
  wire [31:0] w_9 = w_5 ^ w_8; // @[src/main/scala/crypto/aes/KeySchedule.scala 63:21]
  wire [31:0] w_10 = w_6 ^ w_9; // @[src/main/scala/crypto/aes/KeySchedule.scala 63:21]
  wire [31:0] w_11 = w_7 ^ w_10; // @[src/main/scala/crypto/aes/KeySchedule.scala 63:21]
  wire [31:0] _t_T_18 = {w_11[23:0],w_11[31:24]}; // @[src/main/scala/crypto/aes/KeySchedule.scala 23:43]
  wire [7:0] _GEN_2049 = 8'h1 == _t_T_18[15:8] ? 8'h7c : 8'h63; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2050 = 8'h2 == _t_T_18[15:8] ? 8'h77 : _GEN_2049; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2051 = 8'h3 == _t_T_18[15:8] ? 8'h7b : _GEN_2050; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2052 = 8'h4 == _t_T_18[15:8] ? 8'hf2 : _GEN_2051; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2053 = 8'h5 == _t_T_18[15:8] ? 8'h6b : _GEN_2052; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2054 = 8'h6 == _t_T_18[15:8] ? 8'h6f : _GEN_2053; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2055 = 8'h7 == _t_T_18[15:8] ? 8'hc5 : _GEN_2054; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2056 = 8'h8 == _t_T_18[15:8] ? 8'h30 : _GEN_2055; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2057 = 8'h9 == _t_T_18[15:8] ? 8'h1 : _GEN_2056; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2058 = 8'ha == _t_T_18[15:8] ? 8'h67 : _GEN_2057; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2059 = 8'hb == _t_T_18[15:8] ? 8'h2b : _GEN_2058; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2060 = 8'hc == _t_T_18[15:8] ? 8'hfe : _GEN_2059; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2061 = 8'hd == _t_T_18[15:8] ? 8'hd7 : _GEN_2060; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2062 = 8'he == _t_T_18[15:8] ? 8'hab : _GEN_2061; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2063 = 8'hf == _t_T_18[15:8] ? 8'h76 : _GEN_2062; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2064 = 8'h10 == _t_T_18[15:8] ? 8'hca : _GEN_2063; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2065 = 8'h11 == _t_T_18[15:8] ? 8'h82 : _GEN_2064; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2066 = 8'h12 == _t_T_18[15:8] ? 8'hc9 : _GEN_2065; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2067 = 8'h13 == _t_T_18[15:8] ? 8'h7d : _GEN_2066; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2068 = 8'h14 == _t_T_18[15:8] ? 8'hfa : _GEN_2067; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2069 = 8'h15 == _t_T_18[15:8] ? 8'h59 : _GEN_2068; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2070 = 8'h16 == _t_T_18[15:8] ? 8'h47 : _GEN_2069; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2071 = 8'h17 == _t_T_18[15:8] ? 8'hf0 : _GEN_2070; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2072 = 8'h18 == _t_T_18[15:8] ? 8'had : _GEN_2071; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2073 = 8'h19 == _t_T_18[15:8] ? 8'hd4 : _GEN_2072; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2074 = 8'h1a == _t_T_18[15:8] ? 8'ha2 : _GEN_2073; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2075 = 8'h1b == _t_T_18[15:8] ? 8'haf : _GEN_2074; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2076 = 8'h1c == _t_T_18[15:8] ? 8'h9c : _GEN_2075; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2077 = 8'h1d == _t_T_18[15:8] ? 8'ha4 : _GEN_2076; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2078 = 8'h1e == _t_T_18[15:8] ? 8'h72 : _GEN_2077; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2079 = 8'h1f == _t_T_18[15:8] ? 8'hc0 : _GEN_2078; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2080 = 8'h20 == _t_T_18[15:8] ? 8'hb7 : _GEN_2079; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2081 = 8'h21 == _t_T_18[15:8] ? 8'hfd : _GEN_2080; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2082 = 8'h22 == _t_T_18[15:8] ? 8'h93 : _GEN_2081; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2083 = 8'h23 == _t_T_18[15:8] ? 8'h26 : _GEN_2082; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2084 = 8'h24 == _t_T_18[15:8] ? 8'h36 : _GEN_2083; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2085 = 8'h25 == _t_T_18[15:8] ? 8'h3f : _GEN_2084; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2086 = 8'h26 == _t_T_18[15:8] ? 8'hf7 : _GEN_2085; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2087 = 8'h27 == _t_T_18[15:8] ? 8'hcc : _GEN_2086; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2088 = 8'h28 == _t_T_18[15:8] ? 8'h34 : _GEN_2087; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2089 = 8'h29 == _t_T_18[15:8] ? 8'ha5 : _GEN_2088; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2090 = 8'h2a == _t_T_18[15:8] ? 8'he5 : _GEN_2089; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2091 = 8'h2b == _t_T_18[15:8] ? 8'hf1 : _GEN_2090; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2092 = 8'h2c == _t_T_18[15:8] ? 8'h71 : _GEN_2091; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2093 = 8'h2d == _t_T_18[15:8] ? 8'hd8 : _GEN_2092; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2094 = 8'h2e == _t_T_18[15:8] ? 8'h31 : _GEN_2093; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2095 = 8'h2f == _t_T_18[15:8] ? 8'h15 : _GEN_2094; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2096 = 8'h30 == _t_T_18[15:8] ? 8'h4 : _GEN_2095; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2097 = 8'h31 == _t_T_18[15:8] ? 8'hc7 : _GEN_2096; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2098 = 8'h32 == _t_T_18[15:8] ? 8'h23 : _GEN_2097; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2099 = 8'h33 == _t_T_18[15:8] ? 8'hc3 : _GEN_2098; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2100 = 8'h34 == _t_T_18[15:8] ? 8'h18 : _GEN_2099; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2101 = 8'h35 == _t_T_18[15:8] ? 8'h96 : _GEN_2100; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2102 = 8'h36 == _t_T_18[15:8] ? 8'h5 : _GEN_2101; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2103 = 8'h37 == _t_T_18[15:8] ? 8'h9a : _GEN_2102; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2104 = 8'h38 == _t_T_18[15:8] ? 8'h7 : _GEN_2103; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2105 = 8'h39 == _t_T_18[15:8] ? 8'h12 : _GEN_2104; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2106 = 8'h3a == _t_T_18[15:8] ? 8'h80 : _GEN_2105; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2107 = 8'h3b == _t_T_18[15:8] ? 8'he2 : _GEN_2106; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2108 = 8'h3c == _t_T_18[15:8] ? 8'heb : _GEN_2107; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2109 = 8'h3d == _t_T_18[15:8] ? 8'h27 : _GEN_2108; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2110 = 8'h3e == _t_T_18[15:8] ? 8'hb2 : _GEN_2109; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2111 = 8'h3f == _t_T_18[15:8] ? 8'h75 : _GEN_2110; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2112 = 8'h40 == _t_T_18[15:8] ? 8'h9 : _GEN_2111; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2113 = 8'h41 == _t_T_18[15:8] ? 8'h83 : _GEN_2112; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2114 = 8'h42 == _t_T_18[15:8] ? 8'h2c : _GEN_2113; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2115 = 8'h43 == _t_T_18[15:8] ? 8'h1a : _GEN_2114; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2116 = 8'h44 == _t_T_18[15:8] ? 8'h1b : _GEN_2115; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2117 = 8'h45 == _t_T_18[15:8] ? 8'h6e : _GEN_2116; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2118 = 8'h46 == _t_T_18[15:8] ? 8'h5a : _GEN_2117; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2119 = 8'h47 == _t_T_18[15:8] ? 8'ha0 : _GEN_2118; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2120 = 8'h48 == _t_T_18[15:8] ? 8'h52 : _GEN_2119; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2121 = 8'h49 == _t_T_18[15:8] ? 8'h3b : _GEN_2120; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2122 = 8'h4a == _t_T_18[15:8] ? 8'hd6 : _GEN_2121; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2123 = 8'h4b == _t_T_18[15:8] ? 8'hb3 : _GEN_2122; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2124 = 8'h4c == _t_T_18[15:8] ? 8'h29 : _GEN_2123; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2125 = 8'h4d == _t_T_18[15:8] ? 8'he3 : _GEN_2124; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2126 = 8'h4e == _t_T_18[15:8] ? 8'h2f : _GEN_2125; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2127 = 8'h4f == _t_T_18[15:8] ? 8'h84 : _GEN_2126; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2128 = 8'h50 == _t_T_18[15:8] ? 8'h53 : _GEN_2127; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2129 = 8'h51 == _t_T_18[15:8] ? 8'hd1 : _GEN_2128; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2130 = 8'h52 == _t_T_18[15:8] ? 8'h0 : _GEN_2129; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2131 = 8'h53 == _t_T_18[15:8] ? 8'hed : _GEN_2130; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2132 = 8'h54 == _t_T_18[15:8] ? 8'h20 : _GEN_2131; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2133 = 8'h55 == _t_T_18[15:8] ? 8'hfc : _GEN_2132; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2134 = 8'h56 == _t_T_18[15:8] ? 8'hb1 : _GEN_2133; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2135 = 8'h57 == _t_T_18[15:8] ? 8'h5b : _GEN_2134; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2136 = 8'h58 == _t_T_18[15:8] ? 8'h6a : _GEN_2135; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2137 = 8'h59 == _t_T_18[15:8] ? 8'hcb : _GEN_2136; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2138 = 8'h5a == _t_T_18[15:8] ? 8'hbe : _GEN_2137; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2139 = 8'h5b == _t_T_18[15:8] ? 8'h39 : _GEN_2138; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2140 = 8'h5c == _t_T_18[15:8] ? 8'h4a : _GEN_2139; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2141 = 8'h5d == _t_T_18[15:8] ? 8'h4c : _GEN_2140; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2142 = 8'h5e == _t_T_18[15:8] ? 8'h58 : _GEN_2141; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2143 = 8'h5f == _t_T_18[15:8] ? 8'hcf : _GEN_2142; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2144 = 8'h60 == _t_T_18[15:8] ? 8'hd0 : _GEN_2143; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2145 = 8'h61 == _t_T_18[15:8] ? 8'hef : _GEN_2144; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2146 = 8'h62 == _t_T_18[15:8] ? 8'haa : _GEN_2145; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2147 = 8'h63 == _t_T_18[15:8] ? 8'hfb : _GEN_2146; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2148 = 8'h64 == _t_T_18[15:8] ? 8'h43 : _GEN_2147; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2149 = 8'h65 == _t_T_18[15:8] ? 8'h4d : _GEN_2148; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2150 = 8'h66 == _t_T_18[15:8] ? 8'h33 : _GEN_2149; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2151 = 8'h67 == _t_T_18[15:8] ? 8'h85 : _GEN_2150; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2152 = 8'h68 == _t_T_18[15:8] ? 8'h45 : _GEN_2151; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2153 = 8'h69 == _t_T_18[15:8] ? 8'hf9 : _GEN_2152; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2154 = 8'h6a == _t_T_18[15:8] ? 8'h2 : _GEN_2153; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2155 = 8'h6b == _t_T_18[15:8] ? 8'h7f : _GEN_2154; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2156 = 8'h6c == _t_T_18[15:8] ? 8'h50 : _GEN_2155; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2157 = 8'h6d == _t_T_18[15:8] ? 8'h3c : _GEN_2156; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2158 = 8'h6e == _t_T_18[15:8] ? 8'h9f : _GEN_2157; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2159 = 8'h6f == _t_T_18[15:8] ? 8'ha8 : _GEN_2158; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2160 = 8'h70 == _t_T_18[15:8] ? 8'h51 : _GEN_2159; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2161 = 8'h71 == _t_T_18[15:8] ? 8'ha3 : _GEN_2160; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2162 = 8'h72 == _t_T_18[15:8] ? 8'h40 : _GEN_2161; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2163 = 8'h73 == _t_T_18[15:8] ? 8'h8f : _GEN_2162; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2164 = 8'h74 == _t_T_18[15:8] ? 8'h92 : _GEN_2163; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2165 = 8'h75 == _t_T_18[15:8] ? 8'h9d : _GEN_2164; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2166 = 8'h76 == _t_T_18[15:8] ? 8'h38 : _GEN_2165; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2167 = 8'h77 == _t_T_18[15:8] ? 8'hf5 : _GEN_2166; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2168 = 8'h78 == _t_T_18[15:8] ? 8'hbc : _GEN_2167; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2169 = 8'h79 == _t_T_18[15:8] ? 8'hb6 : _GEN_2168; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2170 = 8'h7a == _t_T_18[15:8] ? 8'hda : _GEN_2169; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2171 = 8'h7b == _t_T_18[15:8] ? 8'h21 : _GEN_2170; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2172 = 8'h7c == _t_T_18[15:8] ? 8'h10 : _GEN_2171; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2173 = 8'h7d == _t_T_18[15:8] ? 8'hff : _GEN_2172; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2174 = 8'h7e == _t_T_18[15:8] ? 8'hf3 : _GEN_2173; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2175 = 8'h7f == _t_T_18[15:8] ? 8'hd2 : _GEN_2174; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2176 = 8'h80 == _t_T_18[15:8] ? 8'hcd : _GEN_2175; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2177 = 8'h81 == _t_T_18[15:8] ? 8'hc : _GEN_2176; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2178 = 8'h82 == _t_T_18[15:8] ? 8'h13 : _GEN_2177; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2179 = 8'h83 == _t_T_18[15:8] ? 8'hec : _GEN_2178; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2180 = 8'h84 == _t_T_18[15:8] ? 8'h5f : _GEN_2179; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2181 = 8'h85 == _t_T_18[15:8] ? 8'h97 : _GEN_2180; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2182 = 8'h86 == _t_T_18[15:8] ? 8'h44 : _GEN_2181; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2183 = 8'h87 == _t_T_18[15:8] ? 8'h17 : _GEN_2182; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2184 = 8'h88 == _t_T_18[15:8] ? 8'hc4 : _GEN_2183; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2185 = 8'h89 == _t_T_18[15:8] ? 8'ha7 : _GEN_2184; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2186 = 8'h8a == _t_T_18[15:8] ? 8'h7e : _GEN_2185; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2187 = 8'h8b == _t_T_18[15:8] ? 8'h3d : _GEN_2186; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2188 = 8'h8c == _t_T_18[15:8] ? 8'h64 : _GEN_2187; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2189 = 8'h8d == _t_T_18[15:8] ? 8'h5d : _GEN_2188; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2190 = 8'h8e == _t_T_18[15:8] ? 8'h19 : _GEN_2189; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2191 = 8'h8f == _t_T_18[15:8] ? 8'h73 : _GEN_2190; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2192 = 8'h90 == _t_T_18[15:8] ? 8'h60 : _GEN_2191; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2193 = 8'h91 == _t_T_18[15:8] ? 8'h81 : _GEN_2192; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2194 = 8'h92 == _t_T_18[15:8] ? 8'h4f : _GEN_2193; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2195 = 8'h93 == _t_T_18[15:8] ? 8'hdc : _GEN_2194; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2196 = 8'h94 == _t_T_18[15:8] ? 8'h22 : _GEN_2195; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2197 = 8'h95 == _t_T_18[15:8] ? 8'h2a : _GEN_2196; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2198 = 8'h96 == _t_T_18[15:8] ? 8'h90 : _GEN_2197; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2199 = 8'h97 == _t_T_18[15:8] ? 8'h88 : _GEN_2198; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2200 = 8'h98 == _t_T_18[15:8] ? 8'h46 : _GEN_2199; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2201 = 8'h99 == _t_T_18[15:8] ? 8'hee : _GEN_2200; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2202 = 8'h9a == _t_T_18[15:8] ? 8'hb8 : _GEN_2201; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2203 = 8'h9b == _t_T_18[15:8] ? 8'h14 : _GEN_2202; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2204 = 8'h9c == _t_T_18[15:8] ? 8'hde : _GEN_2203; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2205 = 8'h9d == _t_T_18[15:8] ? 8'h5e : _GEN_2204; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2206 = 8'h9e == _t_T_18[15:8] ? 8'hb : _GEN_2205; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2207 = 8'h9f == _t_T_18[15:8] ? 8'hdb : _GEN_2206; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2208 = 8'ha0 == _t_T_18[15:8] ? 8'he0 : _GEN_2207; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2209 = 8'ha1 == _t_T_18[15:8] ? 8'h32 : _GEN_2208; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2210 = 8'ha2 == _t_T_18[15:8] ? 8'h3a : _GEN_2209; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2211 = 8'ha3 == _t_T_18[15:8] ? 8'ha : _GEN_2210; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2212 = 8'ha4 == _t_T_18[15:8] ? 8'h49 : _GEN_2211; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2213 = 8'ha5 == _t_T_18[15:8] ? 8'h6 : _GEN_2212; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2214 = 8'ha6 == _t_T_18[15:8] ? 8'h24 : _GEN_2213; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2215 = 8'ha7 == _t_T_18[15:8] ? 8'h5c : _GEN_2214; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2216 = 8'ha8 == _t_T_18[15:8] ? 8'hc2 : _GEN_2215; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2217 = 8'ha9 == _t_T_18[15:8] ? 8'hd3 : _GEN_2216; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2218 = 8'haa == _t_T_18[15:8] ? 8'hac : _GEN_2217; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2219 = 8'hab == _t_T_18[15:8] ? 8'h62 : _GEN_2218; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2220 = 8'hac == _t_T_18[15:8] ? 8'h91 : _GEN_2219; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2221 = 8'had == _t_T_18[15:8] ? 8'h95 : _GEN_2220; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2222 = 8'hae == _t_T_18[15:8] ? 8'he4 : _GEN_2221; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2223 = 8'haf == _t_T_18[15:8] ? 8'h79 : _GEN_2222; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2224 = 8'hb0 == _t_T_18[15:8] ? 8'he7 : _GEN_2223; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2225 = 8'hb1 == _t_T_18[15:8] ? 8'hc8 : _GEN_2224; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2226 = 8'hb2 == _t_T_18[15:8] ? 8'h37 : _GEN_2225; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2227 = 8'hb3 == _t_T_18[15:8] ? 8'h6d : _GEN_2226; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2228 = 8'hb4 == _t_T_18[15:8] ? 8'h8d : _GEN_2227; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2229 = 8'hb5 == _t_T_18[15:8] ? 8'hd5 : _GEN_2228; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2230 = 8'hb6 == _t_T_18[15:8] ? 8'h4e : _GEN_2229; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2231 = 8'hb7 == _t_T_18[15:8] ? 8'ha9 : _GEN_2230; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2232 = 8'hb8 == _t_T_18[15:8] ? 8'h6c : _GEN_2231; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2233 = 8'hb9 == _t_T_18[15:8] ? 8'h56 : _GEN_2232; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2234 = 8'hba == _t_T_18[15:8] ? 8'hf4 : _GEN_2233; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2235 = 8'hbb == _t_T_18[15:8] ? 8'hea : _GEN_2234; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2236 = 8'hbc == _t_T_18[15:8] ? 8'h65 : _GEN_2235; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2237 = 8'hbd == _t_T_18[15:8] ? 8'h7a : _GEN_2236; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2238 = 8'hbe == _t_T_18[15:8] ? 8'hae : _GEN_2237; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2239 = 8'hbf == _t_T_18[15:8] ? 8'h8 : _GEN_2238; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2240 = 8'hc0 == _t_T_18[15:8] ? 8'hba : _GEN_2239; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2241 = 8'hc1 == _t_T_18[15:8] ? 8'h78 : _GEN_2240; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2242 = 8'hc2 == _t_T_18[15:8] ? 8'h25 : _GEN_2241; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2243 = 8'hc3 == _t_T_18[15:8] ? 8'h2e : _GEN_2242; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2244 = 8'hc4 == _t_T_18[15:8] ? 8'h1c : _GEN_2243; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2245 = 8'hc5 == _t_T_18[15:8] ? 8'ha6 : _GEN_2244; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2246 = 8'hc6 == _t_T_18[15:8] ? 8'hb4 : _GEN_2245; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2247 = 8'hc7 == _t_T_18[15:8] ? 8'hc6 : _GEN_2246; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2248 = 8'hc8 == _t_T_18[15:8] ? 8'he8 : _GEN_2247; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2249 = 8'hc9 == _t_T_18[15:8] ? 8'hdd : _GEN_2248; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2250 = 8'hca == _t_T_18[15:8] ? 8'h74 : _GEN_2249; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2251 = 8'hcb == _t_T_18[15:8] ? 8'h1f : _GEN_2250; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2252 = 8'hcc == _t_T_18[15:8] ? 8'h4b : _GEN_2251; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2253 = 8'hcd == _t_T_18[15:8] ? 8'hbd : _GEN_2252; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2254 = 8'hce == _t_T_18[15:8] ? 8'h8b : _GEN_2253; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2255 = 8'hcf == _t_T_18[15:8] ? 8'h8a : _GEN_2254; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2256 = 8'hd0 == _t_T_18[15:8] ? 8'h70 : _GEN_2255; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2257 = 8'hd1 == _t_T_18[15:8] ? 8'h3e : _GEN_2256; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2258 = 8'hd2 == _t_T_18[15:8] ? 8'hb5 : _GEN_2257; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2259 = 8'hd3 == _t_T_18[15:8] ? 8'h66 : _GEN_2258; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2260 = 8'hd4 == _t_T_18[15:8] ? 8'h48 : _GEN_2259; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2261 = 8'hd5 == _t_T_18[15:8] ? 8'h3 : _GEN_2260; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2262 = 8'hd6 == _t_T_18[15:8] ? 8'hf6 : _GEN_2261; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2263 = 8'hd7 == _t_T_18[15:8] ? 8'he : _GEN_2262; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2264 = 8'hd8 == _t_T_18[15:8] ? 8'h61 : _GEN_2263; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2265 = 8'hd9 == _t_T_18[15:8] ? 8'h35 : _GEN_2264; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2266 = 8'hda == _t_T_18[15:8] ? 8'h57 : _GEN_2265; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2267 = 8'hdb == _t_T_18[15:8] ? 8'hb9 : _GEN_2266; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2268 = 8'hdc == _t_T_18[15:8] ? 8'h86 : _GEN_2267; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2269 = 8'hdd == _t_T_18[15:8] ? 8'hc1 : _GEN_2268; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2270 = 8'hde == _t_T_18[15:8] ? 8'h1d : _GEN_2269; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2271 = 8'hdf == _t_T_18[15:8] ? 8'h9e : _GEN_2270; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2272 = 8'he0 == _t_T_18[15:8] ? 8'he1 : _GEN_2271; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2273 = 8'he1 == _t_T_18[15:8] ? 8'hf8 : _GEN_2272; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2274 = 8'he2 == _t_T_18[15:8] ? 8'h98 : _GEN_2273; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2275 = 8'he3 == _t_T_18[15:8] ? 8'h11 : _GEN_2274; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2276 = 8'he4 == _t_T_18[15:8] ? 8'h69 : _GEN_2275; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2277 = 8'he5 == _t_T_18[15:8] ? 8'hd9 : _GEN_2276; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2278 = 8'he6 == _t_T_18[15:8] ? 8'h8e : _GEN_2277; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2279 = 8'he7 == _t_T_18[15:8] ? 8'h94 : _GEN_2278; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2280 = 8'he8 == _t_T_18[15:8] ? 8'h9b : _GEN_2279; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2281 = 8'he9 == _t_T_18[15:8] ? 8'h1e : _GEN_2280; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2282 = 8'hea == _t_T_18[15:8] ? 8'h87 : _GEN_2281; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2283 = 8'heb == _t_T_18[15:8] ? 8'he9 : _GEN_2282; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2284 = 8'hec == _t_T_18[15:8] ? 8'hce : _GEN_2283; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2285 = 8'hed == _t_T_18[15:8] ? 8'h55 : _GEN_2284; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2286 = 8'hee == _t_T_18[15:8] ? 8'h28 : _GEN_2285; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2287 = 8'hef == _t_T_18[15:8] ? 8'hdf : _GEN_2286; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2288 = 8'hf0 == _t_T_18[15:8] ? 8'h8c : _GEN_2287; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2289 = 8'hf1 == _t_T_18[15:8] ? 8'ha1 : _GEN_2288; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2290 = 8'hf2 == _t_T_18[15:8] ? 8'h89 : _GEN_2289; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2291 = 8'hf3 == _t_T_18[15:8] ? 8'hd : _GEN_2290; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2292 = 8'hf4 == _t_T_18[15:8] ? 8'hbf : _GEN_2291; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2293 = 8'hf5 == _t_T_18[15:8] ? 8'he6 : _GEN_2292; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2294 = 8'hf6 == _t_T_18[15:8] ? 8'h42 : _GEN_2293; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2295 = 8'hf7 == _t_T_18[15:8] ? 8'h68 : _GEN_2294; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2296 = 8'hf8 == _t_T_18[15:8] ? 8'h41 : _GEN_2295; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2297 = 8'hf9 == _t_T_18[15:8] ? 8'h99 : _GEN_2296; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2298 = 8'hfa == _t_T_18[15:8] ? 8'h2d : _GEN_2297; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2299 = 8'hfb == _t_T_18[15:8] ? 8'hf : _GEN_2298; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2300 = 8'hfc == _t_T_18[15:8] ? 8'hb0 : _GEN_2299; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2301 = 8'hfd == _t_T_18[15:8] ? 8'h54 : _GEN_2300; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2302 = 8'hfe == _t_T_18[15:8] ? 8'hbb : _GEN_2301; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2303 = 8'hff == _t_T_18[15:8] ? 8'h16 : _GEN_2302; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2305 = 8'h1 == _t_T_18[7:0] ? 8'h7c : 8'h63; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2306 = 8'h2 == _t_T_18[7:0] ? 8'h77 : _GEN_2305; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2307 = 8'h3 == _t_T_18[7:0] ? 8'h7b : _GEN_2306; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2308 = 8'h4 == _t_T_18[7:0] ? 8'hf2 : _GEN_2307; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2309 = 8'h5 == _t_T_18[7:0] ? 8'h6b : _GEN_2308; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2310 = 8'h6 == _t_T_18[7:0] ? 8'h6f : _GEN_2309; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2311 = 8'h7 == _t_T_18[7:0] ? 8'hc5 : _GEN_2310; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2312 = 8'h8 == _t_T_18[7:0] ? 8'h30 : _GEN_2311; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2313 = 8'h9 == _t_T_18[7:0] ? 8'h1 : _GEN_2312; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2314 = 8'ha == _t_T_18[7:0] ? 8'h67 : _GEN_2313; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2315 = 8'hb == _t_T_18[7:0] ? 8'h2b : _GEN_2314; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2316 = 8'hc == _t_T_18[7:0] ? 8'hfe : _GEN_2315; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2317 = 8'hd == _t_T_18[7:0] ? 8'hd7 : _GEN_2316; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2318 = 8'he == _t_T_18[7:0] ? 8'hab : _GEN_2317; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2319 = 8'hf == _t_T_18[7:0] ? 8'h76 : _GEN_2318; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2320 = 8'h10 == _t_T_18[7:0] ? 8'hca : _GEN_2319; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2321 = 8'h11 == _t_T_18[7:0] ? 8'h82 : _GEN_2320; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2322 = 8'h12 == _t_T_18[7:0] ? 8'hc9 : _GEN_2321; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2323 = 8'h13 == _t_T_18[7:0] ? 8'h7d : _GEN_2322; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2324 = 8'h14 == _t_T_18[7:0] ? 8'hfa : _GEN_2323; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2325 = 8'h15 == _t_T_18[7:0] ? 8'h59 : _GEN_2324; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2326 = 8'h16 == _t_T_18[7:0] ? 8'h47 : _GEN_2325; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2327 = 8'h17 == _t_T_18[7:0] ? 8'hf0 : _GEN_2326; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2328 = 8'h18 == _t_T_18[7:0] ? 8'had : _GEN_2327; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2329 = 8'h19 == _t_T_18[7:0] ? 8'hd4 : _GEN_2328; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2330 = 8'h1a == _t_T_18[7:0] ? 8'ha2 : _GEN_2329; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2331 = 8'h1b == _t_T_18[7:0] ? 8'haf : _GEN_2330; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2332 = 8'h1c == _t_T_18[7:0] ? 8'h9c : _GEN_2331; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2333 = 8'h1d == _t_T_18[7:0] ? 8'ha4 : _GEN_2332; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2334 = 8'h1e == _t_T_18[7:0] ? 8'h72 : _GEN_2333; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2335 = 8'h1f == _t_T_18[7:0] ? 8'hc0 : _GEN_2334; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2336 = 8'h20 == _t_T_18[7:0] ? 8'hb7 : _GEN_2335; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2337 = 8'h21 == _t_T_18[7:0] ? 8'hfd : _GEN_2336; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2338 = 8'h22 == _t_T_18[7:0] ? 8'h93 : _GEN_2337; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2339 = 8'h23 == _t_T_18[7:0] ? 8'h26 : _GEN_2338; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2340 = 8'h24 == _t_T_18[7:0] ? 8'h36 : _GEN_2339; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2341 = 8'h25 == _t_T_18[7:0] ? 8'h3f : _GEN_2340; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2342 = 8'h26 == _t_T_18[7:0] ? 8'hf7 : _GEN_2341; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2343 = 8'h27 == _t_T_18[7:0] ? 8'hcc : _GEN_2342; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2344 = 8'h28 == _t_T_18[7:0] ? 8'h34 : _GEN_2343; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2345 = 8'h29 == _t_T_18[7:0] ? 8'ha5 : _GEN_2344; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2346 = 8'h2a == _t_T_18[7:0] ? 8'he5 : _GEN_2345; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2347 = 8'h2b == _t_T_18[7:0] ? 8'hf1 : _GEN_2346; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2348 = 8'h2c == _t_T_18[7:0] ? 8'h71 : _GEN_2347; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2349 = 8'h2d == _t_T_18[7:0] ? 8'hd8 : _GEN_2348; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2350 = 8'h2e == _t_T_18[7:0] ? 8'h31 : _GEN_2349; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2351 = 8'h2f == _t_T_18[7:0] ? 8'h15 : _GEN_2350; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2352 = 8'h30 == _t_T_18[7:0] ? 8'h4 : _GEN_2351; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2353 = 8'h31 == _t_T_18[7:0] ? 8'hc7 : _GEN_2352; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2354 = 8'h32 == _t_T_18[7:0] ? 8'h23 : _GEN_2353; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2355 = 8'h33 == _t_T_18[7:0] ? 8'hc3 : _GEN_2354; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2356 = 8'h34 == _t_T_18[7:0] ? 8'h18 : _GEN_2355; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2357 = 8'h35 == _t_T_18[7:0] ? 8'h96 : _GEN_2356; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2358 = 8'h36 == _t_T_18[7:0] ? 8'h5 : _GEN_2357; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2359 = 8'h37 == _t_T_18[7:0] ? 8'h9a : _GEN_2358; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2360 = 8'h38 == _t_T_18[7:0] ? 8'h7 : _GEN_2359; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2361 = 8'h39 == _t_T_18[7:0] ? 8'h12 : _GEN_2360; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2362 = 8'h3a == _t_T_18[7:0] ? 8'h80 : _GEN_2361; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2363 = 8'h3b == _t_T_18[7:0] ? 8'he2 : _GEN_2362; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2364 = 8'h3c == _t_T_18[7:0] ? 8'heb : _GEN_2363; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2365 = 8'h3d == _t_T_18[7:0] ? 8'h27 : _GEN_2364; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2366 = 8'h3e == _t_T_18[7:0] ? 8'hb2 : _GEN_2365; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2367 = 8'h3f == _t_T_18[7:0] ? 8'h75 : _GEN_2366; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2368 = 8'h40 == _t_T_18[7:0] ? 8'h9 : _GEN_2367; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2369 = 8'h41 == _t_T_18[7:0] ? 8'h83 : _GEN_2368; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2370 = 8'h42 == _t_T_18[7:0] ? 8'h2c : _GEN_2369; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2371 = 8'h43 == _t_T_18[7:0] ? 8'h1a : _GEN_2370; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2372 = 8'h44 == _t_T_18[7:0] ? 8'h1b : _GEN_2371; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2373 = 8'h45 == _t_T_18[7:0] ? 8'h6e : _GEN_2372; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2374 = 8'h46 == _t_T_18[7:0] ? 8'h5a : _GEN_2373; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2375 = 8'h47 == _t_T_18[7:0] ? 8'ha0 : _GEN_2374; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2376 = 8'h48 == _t_T_18[7:0] ? 8'h52 : _GEN_2375; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2377 = 8'h49 == _t_T_18[7:0] ? 8'h3b : _GEN_2376; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2378 = 8'h4a == _t_T_18[7:0] ? 8'hd6 : _GEN_2377; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2379 = 8'h4b == _t_T_18[7:0] ? 8'hb3 : _GEN_2378; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2380 = 8'h4c == _t_T_18[7:0] ? 8'h29 : _GEN_2379; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2381 = 8'h4d == _t_T_18[7:0] ? 8'he3 : _GEN_2380; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2382 = 8'h4e == _t_T_18[7:0] ? 8'h2f : _GEN_2381; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2383 = 8'h4f == _t_T_18[7:0] ? 8'h84 : _GEN_2382; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2384 = 8'h50 == _t_T_18[7:0] ? 8'h53 : _GEN_2383; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2385 = 8'h51 == _t_T_18[7:0] ? 8'hd1 : _GEN_2384; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2386 = 8'h52 == _t_T_18[7:0] ? 8'h0 : _GEN_2385; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2387 = 8'h53 == _t_T_18[7:0] ? 8'hed : _GEN_2386; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2388 = 8'h54 == _t_T_18[7:0] ? 8'h20 : _GEN_2387; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2389 = 8'h55 == _t_T_18[7:0] ? 8'hfc : _GEN_2388; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2390 = 8'h56 == _t_T_18[7:0] ? 8'hb1 : _GEN_2389; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2391 = 8'h57 == _t_T_18[7:0] ? 8'h5b : _GEN_2390; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2392 = 8'h58 == _t_T_18[7:0] ? 8'h6a : _GEN_2391; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2393 = 8'h59 == _t_T_18[7:0] ? 8'hcb : _GEN_2392; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2394 = 8'h5a == _t_T_18[7:0] ? 8'hbe : _GEN_2393; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2395 = 8'h5b == _t_T_18[7:0] ? 8'h39 : _GEN_2394; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2396 = 8'h5c == _t_T_18[7:0] ? 8'h4a : _GEN_2395; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2397 = 8'h5d == _t_T_18[7:0] ? 8'h4c : _GEN_2396; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2398 = 8'h5e == _t_T_18[7:0] ? 8'h58 : _GEN_2397; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2399 = 8'h5f == _t_T_18[7:0] ? 8'hcf : _GEN_2398; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2400 = 8'h60 == _t_T_18[7:0] ? 8'hd0 : _GEN_2399; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2401 = 8'h61 == _t_T_18[7:0] ? 8'hef : _GEN_2400; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2402 = 8'h62 == _t_T_18[7:0] ? 8'haa : _GEN_2401; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2403 = 8'h63 == _t_T_18[7:0] ? 8'hfb : _GEN_2402; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2404 = 8'h64 == _t_T_18[7:0] ? 8'h43 : _GEN_2403; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2405 = 8'h65 == _t_T_18[7:0] ? 8'h4d : _GEN_2404; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2406 = 8'h66 == _t_T_18[7:0] ? 8'h33 : _GEN_2405; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2407 = 8'h67 == _t_T_18[7:0] ? 8'h85 : _GEN_2406; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2408 = 8'h68 == _t_T_18[7:0] ? 8'h45 : _GEN_2407; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2409 = 8'h69 == _t_T_18[7:0] ? 8'hf9 : _GEN_2408; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2410 = 8'h6a == _t_T_18[7:0] ? 8'h2 : _GEN_2409; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2411 = 8'h6b == _t_T_18[7:0] ? 8'h7f : _GEN_2410; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2412 = 8'h6c == _t_T_18[7:0] ? 8'h50 : _GEN_2411; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2413 = 8'h6d == _t_T_18[7:0] ? 8'h3c : _GEN_2412; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2414 = 8'h6e == _t_T_18[7:0] ? 8'h9f : _GEN_2413; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2415 = 8'h6f == _t_T_18[7:0] ? 8'ha8 : _GEN_2414; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2416 = 8'h70 == _t_T_18[7:0] ? 8'h51 : _GEN_2415; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2417 = 8'h71 == _t_T_18[7:0] ? 8'ha3 : _GEN_2416; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2418 = 8'h72 == _t_T_18[7:0] ? 8'h40 : _GEN_2417; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2419 = 8'h73 == _t_T_18[7:0] ? 8'h8f : _GEN_2418; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2420 = 8'h74 == _t_T_18[7:0] ? 8'h92 : _GEN_2419; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2421 = 8'h75 == _t_T_18[7:0] ? 8'h9d : _GEN_2420; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2422 = 8'h76 == _t_T_18[7:0] ? 8'h38 : _GEN_2421; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2423 = 8'h77 == _t_T_18[7:0] ? 8'hf5 : _GEN_2422; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2424 = 8'h78 == _t_T_18[7:0] ? 8'hbc : _GEN_2423; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2425 = 8'h79 == _t_T_18[7:0] ? 8'hb6 : _GEN_2424; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2426 = 8'h7a == _t_T_18[7:0] ? 8'hda : _GEN_2425; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2427 = 8'h7b == _t_T_18[7:0] ? 8'h21 : _GEN_2426; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2428 = 8'h7c == _t_T_18[7:0] ? 8'h10 : _GEN_2427; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2429 = 8'h7d == _t_T_18[7:0] ? 8'hff : _GEN_2428; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2430 = 8'h7e == _t_T_18[7:0] ? 8'hf3 : _GEN_2429; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2431 = 8'h7f == _t_T_18[7:0] ? 8'hd2 : _GEN_2430; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2432 = 8'h80 == _t_T_18[7:0] ? 8'hcd : _GEN_2431; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2433 = 8'h81 == _t_T_18[7:0] ? 8'hc : _GEN_2432; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2434 = 8'h82 == _t_T_18[7:0] ? 8'h13 : _GEN_2433; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2435 = 8'h83 == _t_T_18[7:0] ? 8'hec : _GEN_2434; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2436 = 8'h84 == _t_T_18[7:0] ? 8'h5f : _GEN_2435; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2437 = 8'h85 == _t_T_18[7:0] ? 8'h97 : _GEN_2436; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2438 = 8'h86 == _t_T_18[7:0] ? 8'h44 : _GEN_2437; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2439 = 8'h87 == _t_T_18[7:0] ? 8'h17 : _GEN_2438; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2440 = 8'h88 == _t_T_18[7:0] ? 8'hc4 : _GEN_2439; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2441 = 8'h89 == _t_T_18[7:0] ? 8'ha7 : _GEN_2440; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2442 = 8'h8a == _t_T_18[7:0] ? 8'h7e : _GEN_2441; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2443 = 8'h8b == _t_T_18[7:0] ? 8'h3d : _GEN_2442; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2444 = 8'h8c == _t_T_18[7:0] ? 8'h64 : _GEN_2443; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2445 = 8'h8d == _t_T_18[7:0] ? 8'h5d : _GEN_2444; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2446 = 8'h8e == _t_T_18[7:0] ? 8'h19 : _GEN_2445; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2447 = 8'h8f == _t_T_18[7:0] ? 8'h73 : _GEN_2446; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2448 = 8'h90 == _t_T_18[7:0] ? 8'h60 : _GEN_2447; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2449 = 8'h91 == _t_T_18[7:0] ? 8'h81 : _GEN_2448; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2450 = 8'h92 == _t_T_18[7:0] ? 8'h4f : _GEN_2449; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2451 = 8'h93 == _t_T_18[7:0] ? 8'hdc : _GEN_2450; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2452 = 8'h94 == _t_T_18[7:0] ? 8'h22 : _GEN_2451; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2453 = 8'h95 == _t_T_18[7:0] ? 8'h2a : _GEN_2452; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2454 = 8'h96 == _t_T_18[7:0] ? 8'h90 : _GEN_2453; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2455 = 8'h97 == _t_T_18[7:0] ? 8'h88 : _GEN_2454; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2456 = 8'h98 == _t_T_18[7:0] ? 8'h46 : _GEN_2455; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2457 = 8'h99 == _t_T_18[7:0] ? 8'hee : _GEN_2456; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2458 = 8'h9a == _t_T_18[7:0] ? 8'hb8 : _GEN_2457; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2459 = 8'h9b == _t_T_18[7:0] ? 8'h14 : _GEN_2458; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2460 = 8'h9c == _t_T_18[7:0] ? 8'hde : _GEN_2459; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2461 = 8'h9d == _t_T_18[7:0] ? 8'h5e : _GEN_2460; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2462 = 8'h9e == _t_T_18[7:0] ? 8'hb : _GEN_2461; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2463 = 8'h9f == _t_T_18[7:0] ? 8'hdb : _GEN_2462; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2464 = 8'ha0 == _t_T_18[7:0] ? 8'he0 : _GEN_2463; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2465 = 8'ha1 == _t_T_18[7:0] ? 8'h32 : _GEN_2464; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2466 = 8'ha2 == _t_T_18[7:0] ? 8'h3a : _GEN_2465; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2467 = 8'ha3 == _t_T_18[7:0] ? 8'ha : _GEN_2466; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2468 = 8'ha4 == _t_T_18[7:0] ? 8'h49 : _GEN_2467; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2469 = 8'ha5 == _t_T_18[7:0] ? 8'h6 : _GEN_2468; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2470 = 8'ha6 == _t_T_18[7:0] ? 8'h24 : _GEN_2469; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2471 = 8'ha7 == _t_T_18[7:0] ? 8'h5c : _GEN_2470; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2472 = 8'ha8 == _t_T_18[7:0] ? 8'hc2 : _GEN_2471; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2473 = 8'ha9 == _t_T_18[7:0] ? 8'hd3 : _GEN_2472; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2474 = 8'haa == _t_T_18[7:0] ? 8'hac : _GEN_2473; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2475 = 8'hab == _t_T_18[7:0] ? 8'h62 : _GEN_2474; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2476 = 8'hac == _t_T_18[7:0] ? 8'h91 : _GEN_2475; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2477 = 8'had == _t_T_18[7:0] ? 8'h95 : _GEN_2476; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2478 = 8'hae == _t_T_18[7:0] ? 8'he4 : _GEN_2477; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2479 = 8'haf == _t_T_18[7:0] ? 8'h79 : _GEN_2478; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2480 = 8'hb0 == _t_T_18[7:0] ? 8'he7 : _GEN_2479; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2481 = 8'hb1 == _t_T_18[7:0] ? 8'hc8 : _GEN_2480; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2482 = 8'hb2 == _t_T_18[7:0] ? 8'h37 : _GEN_2481; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2483 = 8'hb3 == _t_T_18[7:0] ? 8'h6d : _GEN_2482; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2484 = 8'hb4 == _t_T_18[7:0] ? 8'h8d : _GEN_2483; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2485 = 8'hb5 == _t_T_18[7:0] ? 8'hd5 : _GEN_2484; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2486 = 8'hb6 == _t_T_18[7:0] ? 8'h4e : _GEN_2485; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2487 = 8'hb7 == _t_T_18[7:0] ? 8'ha9 : _GEN_2486; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2488 = 8'hb8 == _t_T_18[7:0] ? 8'h6c : _GEN_2487; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2489 = 8'hb9 == _t_T_18[7:0] ? 8'h56 : _GEN_2488; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2490 = 8'hba == _t_T_18[7:0] ? 8'hf4 : _GEN_2489; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2491 = 8'hbb == _t_T_18[7:0] ? 8'hea : _GEN_2490; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2492 = 8'hbc == _t_T_18[7:0] ? 8'h65 : _GEN_2491; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2493 = 8'hbd == _t_T_18[7:0] ? 8'h7a : _GEN_2492; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2494 = 8'hbe == _t_T_18[7:0] ? 8'hae : _GEN_2493; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2495 = 8'hbf == _t_T_18[7:0] ? 8'h8 : _GEN_2494; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2496 = 8'hc0 == _t_T_18[7:0] ? 8'hba : _GEN_2495; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2497 = 8'hc1 == _t_T_18[7:0] ? 8'h78 : _GEN_2496; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2498 = 8'hc2 == _t_T_18[7:0] ? 8'h25 : _GEN_2497; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2499 = 8'hc3 == _t_T_18[7:0] ? 8'h2e : _GEN_2498; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2500 = 8'hc4 == _t_T_18[7:0] ? 8'h1c : _GEN_2499; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2501 = 8'hc5 == _t_T_18[7:0] ? 8'ha6 : _GEN_2500; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2502 = 8'hc6 == _t_T_18[7:0] ? 8'hb4 : _GEN_2501; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2503 = 8'hc7 == _t_T_18[7:0] ? 8'hc6 : _GEN_2502; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2504 = 8'hc8 == _t_T_18[7:0] ? 8'he8 : _GEN_2503; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2505 = 8'hc9 == _t_T_18[7:0] ? 8'hdd : _GEN_2504; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2506 = 8'hca == _t_T_18[7:0] ? 8'h74 : _GEN_2505; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2507 = 8'hcb == _t_T_18[7:0] ? 8'h1f : _GEN_2506; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2508 = 8'hcc == _t_T_18[7:0] ? 8'h4b : _GEN_2507; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2509 = 8'hcd == _t_T_18[7:0] ? 8'hbd : _GEN_2508; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2510 = 8'hce == _t_T_18[7:0] ? 8'h8b : _GEN_2509; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2511 = 8'hcf == _t_T_18[7:0] ? 8'h8a : _GEN_2510; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2512 = 8'hd0 == _t_T_18[7:0] ? 8'h70 : _GEN_2511; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2513 = 8'hd1 == _t_T_18[7:0] ? 8'h3e : _GEN_2512; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2514 = 8'hd2 == _t_T_18[7:0] ? 8'hb5 : _GEN_2513; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2515 = 8'hd3 == _t_T_18[7:0] ? 8'h66 : _GEN_2514; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2516 = 8'hd4 == _t_T_18[7:0] ? 8'h48 : _GEN_2515; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2517 = 8'hd5 == _t_T_18[7:0] ? 8'h3 : _GEN_2516; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2518 = 8'hd6 == _t_T_18[7:0] ? 8'hf6 : _GEN_2517; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2519 = 8'hd7 == _t_T_18[7:0] ? 8'he : _GEN_2518; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2520 = 8'hd8 == _t_T_18[7:0] ? 8'h61 : _GEN_2519; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2521 = 8'hd9 == _t_T_18[7:0] ? 8'h35 : _GEN_2520; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2522 = 8'hda == _t_T_18[7:0] ? 8'h57 : _GEN_2521; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2523 = 8'hdb == _t_T_18[7:0] ? 8'hb9 : _GEN_2522; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2524 = 8'hdc == _t_T_18[7:0] ? 8'h86 : _GEN_2523; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2525 = 8'hdd == _t_T_18[7:0] ? 8'hc1 : _GEN_2524; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2526 = 8'hde == _t_T_18[7:0] ? 8'h1d : _GEN_2525; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2527 = 8'hdf == _t_T_18[7:0] ? 8'h9e : _GEN_2526; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2528 = 8'he0 == _t_T_18[7:0] ? 8'he1 : _GEN_2527; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2529 = 8'he1 == _t_T_18[7:0] ? 8'hf8 : _GEN_2528; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2530 = 8'he2 == _t_T_18[7:0] ? 8'h98 : _GEN_2529; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2531 = 8'he3 == _t_T_18[7:0] ? 8'h11 : _GEN_2530; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2532 = 8'he4 == _t_T_18[7:0] ? 8'h69 : _GEN_2531; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2533 = 8'he5 == _t_T_18[7:0] ? 8'hd9 : _GEN_2532; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2534 = 8'he6 == _t_T_18[7:0] ? 8'h8e : _GEN_2533; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2535 = 8'he7 == _t_T_18[7:0] ? 8'h94 : _GEN_2534; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2536 = 8'he8 == _t_T_18[7:0] ? 8'h9b : _GEN_2535; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2537 = 8'he9 == _t_T_18[7:0] ? 8'h1e : _GEN_2536; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2538 = 8'hea == _t_T_18[7:0] ? 8'h87 : _GEN_2537; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2539 = 8'heb == _t_T_18[7:0] ? 8'he9 : _GEN_2538; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2540 = 8'hec == _t_T_18[7:0] ? 8'hce : _GEN_2539; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2541 = 8'hed == _t_T_18[7:0] ? 8'h55 : _GEN_2540; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2542 = 8'hee == _t_T_18[7:0] ? 8'h28 : _GEN_2541; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2543 = 8'hef == _t_T_18[7:0] ? 8'hdf : _GEN_2542; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2544 = 8'hf0 == _t_T_18[7:0] ? 8'h8c : _GEN_2543; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2545 = 8'hf1 == _t_T_18[7:0] ? 8'ha1 : _GEN_2544; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2546 = 8'hf2 == _t_T_18[7:0] ? 8'h89 : _GEN_2545; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2547 = 8'hf3 == _t_T_18[7:0] ? 8'hd : _GEN_2546; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2548 = 8'hf4 == _t_T_18[7:0] ? 8'hbf : _GEN_2547; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2549 = 8'hf5 == _t_T_18[7:0] ? 8'he6 : _GEN_2548; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2550 = 8'hf6 == _t_T_18[7:0] ? 8'h42 : _GEN_2549; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2551 = 8'hf7 == _t_T_18[7:0] ? 8'h68 : _GEN_2550; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2552 = 8'hf8 == _t_T_18[7:0] ? 8'h41 : _GEN_2551; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2553 = 8'hf9 == _t_T_18[7:0] ? 8'h99 : _GEN_2552; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2554 = 8'hfa == _t_T_18[7:0] ? 8'h2d : _GEN_2553; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2555 = 8'hfb == _t_T_18[7:0] ? 8'hf : _GEN_2554; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2556 = 8'hfc == _t_T_18[7:0] ? 8'hb0 : _GEN_2555; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2557 = 8'hfd == _t_T_18[7:0] ? 8'h54 : _GEN_2556; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2558 = 8'hfe == _t_T_18[7:0] ? 8'hbb : _GEN_2557; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2559 = 8'hff == _t_T_18[7:0] ? 8'h16 : _GEN_2558; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2561 = 8'h1 == _t_T_18[31:24] ? 8'h7c : 8'h63; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2562 = 8'h2 == _t_T_18[31:24] ? 8'h77 : _GEN_2561; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2563 = 8'h3 == _t_T_18[31:24] ? 8'h7b : _GEN_2562; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2564 = 8'h4 == _t_T_18[31:24] ? 8'hf2 : _GEN_2563; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2565 = 8'h5 == _t_T_18[31:24] ? 8'h6b : _GEN_2564; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2566 = 8'h6 == _t_T_18[31:24] ? 8'h6f : _GEN_2565; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2567 = 8'h7 == _t_T_18[31:24] ? 8'hc5 : _GEN_2566; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2568 = 8'h8 == _t_T_18[31:24] ? 8'h30 : _GEN_2567; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2569 = 8'h9 == _t_T_18[31:24] ? 8'h1 : _GEN_2568; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2570 = 8'ha == _t_T_18[31:24] ? 8'h67 : _GEN_2569; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2571 = 8'hb == _t_T_18[31:24] ? 8'h2b : _GEN_2570; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2572 = 8'hc == _t_T_18[31:24] ? 8'hfe : _GEN_2571; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2573 = 8'hd == _t_T_18[31:24] ? 8'hd7 : _GEN_2572; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2574 = 8'he == _t_T_18[31:24] ? 8'hab : _GEN_2573; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2575 = 8'hf == _t_T_18[31:24] ? 8'h76 : _GEN_2574; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2576 = 8'h10 == _t_T_18[31:24] ? 8'hca : _GEN_2575; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2577 = 8'h11 == _t_T_18[31:24] ? 8'h82 : _GEN_2576; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2578 = 8'h12 == _t_T_18[31:24] ? 8'hc9 : _GEN_2577; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2579 = 8'h13 == _t_T_18[31:24] ? 8'h7d : _GEN_2578; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2580 = 8'h14 == _t_T_18[31:24] ? 8'hfa : _GEN_2579; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2581 = 8'h15 == _t_T_18[31:24] ? 8'h59 : _GEN_2580; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2582 = 8'h16 == _t_T_18[31:24] ? 8'h47 : _GEN_2581; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2583 = 8'h17 == _t_T_18[31:24] ? 8'hf0 : _GEN_2582; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2584 = 8'h18 == _t_T_18[31:24] ? 8'had : _GEN_2583; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2585 = 8'h19 == _t_T_18[31:24] ? 8'hd4 : _GEN_2584; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2586 = 8'h1a == _t_T_18[31:24] ? 8'ha2 : _GEN_2585; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2587 = 8'h1b == _t_T_18[31:24] ? 8'haf : _GEN_2586; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2588 = 8'h1c == _t_T_18[31:24] ? 8'h9c : _GEN_2587; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2589 = 8'h1d == _t_T_18[31:24] ? 8'ha4 : _GEN_2588; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2590 = 8'h1e == _t_T_18[31:24] ? 8'h72 : _GEN_2589; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2591 = 8'h1f == _t_T_18[31:24] ? 8'hc0 : _GEN_2590; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2592 = 8'h20 == _t_T_18[31:24] ? 8'hb7 : _GEN_2591; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2593 = 8'h21 == _t_T_18[31:24] ? 8'hfd : _GEN_2592; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2594 = 8'h22 == _t_T_18[31:24] ? 8'h93 : _GEN_2593; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2595 = 8'h23 == _t_T_18[31:24] ? 8'h26 : _GEN_2594; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2596 = 8'h24 == _t_T_18[31:24] ? 8'h36 : _GEN_2595; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2597 = 8'h25 == _t_T_18[31:24] ? 8'h3f : _GEN_2596; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2598 = 8'h26 == _t_T_18[31:24] ? 8'hf7 : _GEN_2597; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2599 = 8'h27 == _t_T_18[31:24] ? 8'hcc : _GEN_2598; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2600 = 8'h28 == _t_T_18[31:24] ? 8'h34 : _GEN_2599; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2601 = 8'h29 == _t_T_18[31:24] ? 8'ha5 : _GEN_2600; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2602 = 8'h2a == _t_T_18[31:24] ? 8'he5 : _GEN_2601; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2603 = 8'h2b == _t_T_18[31:24] ? 8'hf1 : _GEN_2602; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2604 = 8'h2c == _t_T_18[31:24] ? 8'h71 : _GEN_2603; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2605 = 8'h2d == _t_T_18[31:24] ? 8'hd8 : _GEN_2604; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2606 = 8'h2e == _t_T_18[31:24] ? 8'h31 : _GEN_2605; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2607 = 8'h2f == _t_T_18[31:24] ? 8'h15 : _GEN_2606; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2608 = 8'h30 == _t_T_18[31:24] ? 8'h4 : _GEN_2607; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2609 = 8'h31 == _t_T_18[31:24] ? 8'hc7 : _GEN_2608; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2610 = 8'h32 == _t_T_18[31:24] ? 8'h23 : _GEN_2609; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2611 = 8'h33 == _t_T_18[31:24] ? 8'hc3 : _GEN_2610; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2612 = 8'h34 == _t_T_18[31:24] ? 8'h18 : _GEN_2611; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2613 = 8'h35 == _t_T_18[31:24] ? 8'h96 : _GEN_2612; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2614 = 8'h36 == _t_T_18[31:24] ? 8'h5 : _GEN_2613; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2615 = 8'h37 == _t_T_18[31:24] ? 8'h9a : _GEN_2614; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2616 = 8'h38 == _t_T_18[31:24] ? 8'h7 : _GEN_2615; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2617 = 8'h39 == _t_T_18[31:24] ? 8'h12 : _GEN_2616; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2618 = 8'h3a == _t_T_18[31:24] ? 8'h80 : _GEN_2617; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2619 = 8'h3b == _t_T_18[31:24] ? 8'he2 : _GEN_2618; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2620 = 8'h3c == _t_T_18[31:24] ? 8'heb : _GEN_2619; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2621 = 8'h3d == _t_T_18[31:24] ? 8'h27 : _GEN_2620; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2622 = 8'h3e == _t_T_18[31:24] ? 8'hb2 : _GEN_2621; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2623 = 8'h3f == _t_T_18[31:24] ? 8'h75 : _GEN_2622; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2624 = 8'h40 == _t_T_18[31:24] ? 8'h9 : _GEN_2623; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2625 = 8'h41 == _t_T_18[31:24] ? 8'h83 : _GEN_2624; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2626 = 8'h42 == _t_T_18[31:24] ? 8'h2c : _GEN_2625; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2627 = 8'h43 == _t_T_18[31:24] ? 8'h1a : _GEN_2626; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2628 = 8'h44 == _t_T_18[31:24] ? 8'h1b : _GEN_2627; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2629 = 8'h45 == _t_T_18[31:24] ? 8'h6e : _GEN_2628; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2630 = 8'h46 == _t_T_18[31:24] ? 8'h5a : _GEN_2629; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2631 = 8'h47 == _t_T_18[31:24] ? 8'ha0 : _GEN_2630; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2632 = 8'h48 == _t_T_18[31:24] ? 8'h52 : _GEN_2631; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2633 = 8'h49 == _t_T_18[31:24] ? 8'h3b : _GEN_2632; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2634 = 8'h4a == _t_T_18[31:24] ? 8'hd6 : _GEN_2633; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2635 = 8'h4b == _t_T_18[31:24] ? 8'hb3 : _GEN_2634; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2636 = 8'h4c == _t_T_18[31:24] ? 8'h29 : _GEN_2635; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2637 = 8'h4d == _t_T_18[31:24] ? 8'he3 : _GEN_2636; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2638 = 8'h4e == _t_T_18[31:24] ? 8'h2f : _GEN_2637; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2639 = 8'h4f == _t_T_18[31:24] ? 8'h84 : _GEN_2638; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2640 = 8'h50 == _t_T_18[31:24] ? 8'h53 : _GEN_2639; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2641 = 8'h51 == _t_T_18[31:24] ? 8'hd1 : _GEN_2640; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2642 = 8'h52 == _t_T_18[31:24] ? 8'h0 : _GEN_2641; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2643 = 8'h53 == _t_T_18[31:24] ? 8'hed : _GEN_2642; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2644 = 8'h54 == _t_T_18[31:24] ? 8'h20 : _GEN_2643; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2645 = 8'h55 == _t_T_18[31:24] ? 8'hfc : _GEN_2644; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2646 = 8'h56 == _t_T_18[31:24] ? 8'hb1 : _GEN_2645; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2647 = 8'h57 == _t_T_18[31:24] ? 8'h5b : _GEN_2646; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2648 = 8'h58 == _t_T_18[31:24] ? 8'h6a : _GEN_2647; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2649 = 8'h59 == _t_T_18[31:24] ? 8'hcb : _GEN_2648; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2650 = 8'h5a == _t_T_18[31:24] ? 8'hbe : _GEN_2649; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2651 = 8'h5b == _t_T_18[31:24] ? 8'h39 : _GEN_2650; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2652 = 8'h5c == _t_T_18[31:24] ? 8'h4a : _GEN_2651; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2653 = 8'h5d == _t_T_18[31:24] ? 8'h4c : _GEN_2652; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2654 = 8'h5e == _t_T_18[31:24] ? 8'h58 : _GEN_2653; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2655 = 8'h5f == _t_T_18[31:24] ? 8'hcf : _GEN_2654; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2656 = 8'h60 == _t_T_18[31:24] ? 8'hd0 : _GEN_2655; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2657 = 8'h61 == _t_T_18[31:24] ? 8'hef : _GEN_2656; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2658 = 8'h62 == _t_T_18[31:24] ? 8'haa : _GEN_2657; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2659 = 8'h63 == _t_T_18[31:24] ? 8'hfb : _GEN_2658; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2660 = 8'h64 == _t_T_18[31:24] ? 8'h43 : _GEN_2659; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2661 = 8'h65 == _t_T_18[31:24] ? 8'h4d : _GEN_2660; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2662 = 8'h66 == _t_T_18[31:24] ? 8'h33 : _GEN_2661; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2663 = 8'h67 == _t_T_18[31:24] ? 8'h85 : _GEN_2662; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2664 = 8'h68 == _t_T_18[31:24] ? 8'h45 : _GEN_2663; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2665 = 8'h69 == _t_T_18[31:24] ? 8'hf9 : _GEN_2664; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2666 = 8'h6a == _t_T_18[31:24] ? 8'h2 : _GEN_2665; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2667 = 8'h6b == _t_T_18[31:24] ? 8'h7f : _GEN_2666; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2668 = 8'h6c == _t_T_18[31:24] ? 8'h50 : _GEN_2667; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2669 = 8'h6d == _t_T_18[31:24] ? 8'h3c : _GEN_2668; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2670 = 8'h6e == _t_T_18[31:24] ? 8'h9f : _GEN_2669; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2671 = 8'h6f == _t_T_18[31:24] ? 8'ha8 : _GEN_2670; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2672 = 8'h70 == _t_T_18[31:24] ? 8'h51 : _GEN_2671; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2673 = 8'h71 == _t_T_18[31:24] ? 8'ha3 : _GEN_2672; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2674 = 8'h72 == _t_T_18[31:24] ? 8'h40 : _GEN_2673; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2675 = 8'h73 == _t_T_18[31:24] ? 8'h8f : _GEN_2674; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2676 = 8'h74 == _t_T_18[31:24] ? 8'h92 : _GEN_2675; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2677 = 8'h75 == _t_T_18[31:24] ? 8'h9d : _GEN_2676; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2678 = 8'h76 == _t_T_18[31:24] ? 8'h38 : _GEN_2677; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2679 = 8'h77 == _t_T_18[31:24] ? 8'hf5 : _GEN_2678; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2680 = 8'h78 == _t_T_18[31:24] ? 8'hbc : _GEN_2679; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2681 = 8'h79 == _t_T_18[31:24] ? 8'hb6 : _GEN_2680; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2682 = 8'h7a == _t_T_18[31:24] ? 8'hda : _GEN_2681; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2683 = 8'h7b == _t_T_18[31:24] ? 8'h21 : _GEN_2682; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2684 = 8'h7c == _t_T_18[31:24] ? 8'h10 : _GEN_2683; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2685 = 8'h7d == _t_T_18[31:24] ? 8'hff : _GEN_2684; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2686 = 8'h7e == _t_T_18[31:24] ? 8'hf3 : _GEN_2685; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2687 = 8'h7f == _t_T_18[31:24] ? 8'hd2 : _GEN_2686; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2688 = 8'h80 == _t_T_18[31:24] ? 8'hcd : _GEN_2687; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2689 = 8'h81 == _t_T_18[31:24] ? 8'hc : _GEN_2688; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2690 = 8'h82 == _t_T_18[31:24] ? 8'h13 : _GEN_2689; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2691 = 8'h83 == _t_T_18[31:24] ? 8'hec : _GEN_2690; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2692 = 8'h84 == _t_T_18[31:24] ? 8'h5f : _GEN_2691; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2693 = 8'h85 == _t_T_18[31:24] ? 8'h97 : _GEN_2692; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2694 = 8'h86 == _t_T_18[31:24] ? 8'h44 : _GEN_2693; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2695 = 8'h87 == _t_T_18[31:24] ? 8'h17 : _GEN_2694; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2696 = 8'h88 == _t_T_18[31:24] ? 8'hc4 : _GEN_2695; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2697 = 8'h89 == _t_T_18[31:24] ? 8'ha7 : _GEN_2696; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2698 = 8'h8a == _t_T_18[31:24] ? 8'h7e : _GEN_2697; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2699 = 8'h8b == _t_T_18[31:24] ? 8'h3d : _GEN_2698; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2700 = 8'h8c == _t_T_18[31:24] ? 8'h64 : _GEN_2699; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2701 = 8'h8d == _t_T_18[31:24] ? 8'h5d : _GEN_2700; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2702 = 8'h8e == _t_T_18[31:24] ? 8'h19 : _GEN_2701; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2703 = 8'h8f == _t_T_18[31:24] ? 8'h73 : _GEN_2702; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2704 = 8'h90 == _t_T_18[31:24] ? 8'h60 : _GEN_2703; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2705 = 8'h91 == _t_T_18[31:24] ? 8'h81 : _GEN_2704; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2706 = 8'h92 == _t_T_18[31:24] ? 8'h4f : _GEN_2705; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2707 = 8'h93 == _t_T_18[31:24] ? 8'hdc : _GEN_2706; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2708 = 8'h94 == _t_T_18[31:24] ? 8'h22 : _GEN_2707; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2709 = 8'h95 == _t_T_18[31:24] ? 8'h2a : _GEN_2708; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2710 = 8'h96 == _t_T_18[31:24] ? 8'h90 : _GEN_2709; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2711 = 8'h97 == _t_T_18[31:24] ? 8'h88 : _GEN_2710; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2712 = 8'h98 == _t_T_18[31:24] ? 8'h46 : _GEN_2711; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2713 = 8'h99 == _t_T_18[31:24] ? 8'hee : _GEN_2712; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2714 = 8'h9a == _t_T_18[31:24] ? 8'hb8 : _GEN_2713; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2715 = 8'h9b == _t_T_18[31:24] ? 8'h14 : _GEN_2714; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2716 = 8'h9c == _t_T_18[31:24] ? 8'hde : _GEN_2715; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2717 = 8'h9d == _t_T_18[31:24] ? 8'h5e : _GEN_2716; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2718 = 8'h9e == _t_T_18[31:24] ? 8'hb : _GEN_2717; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2719 = 8'h9f == _t_T_18[31:24] ? 8'hdb : _GEN_2718; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2720 = 8'ha0 == _t_T_18[31:24] ? 8'he0 : _GEN_2719; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2721 = 8'ha1 == _t_T_18[31:24] ? 8'h32 : _GEN_2720; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2722 = 8'ha2 == _t_T_18[31:24] ? 8'h3a : _GEN_2721; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2723 = 8'ha3 == _t_T_18[31:24] ? 8'ha : _GEN_2722; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2724 = 8'ha4 == _t_T_18[31:24] ? 8'h49 : _GEN_2723; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2725 = 8'ha5 == _t_T_18[31:24] ? 8'h6 : _GEN_2724; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2726 = 8'ha6 == _t_T_18[31:24] ? 8'h24 : _GEN_2725; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2727 = 8'ha7 == _t_T_18[31:24] ? 8'h5c : _GEN_2726; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2728 = 8'ha8 == _t_T_18[31:24] ? 8'hc2 : _GEN_2727; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2729 = 8'ha9 == _t_T_18[31:24] ? 8'hd3 : _GEN_2728; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2730 = 8'haa == _t_T_18[31:24] ? 8'hac : _GEN_2729; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2731 = 8'hab == _t_T_18[31:24] ? 8'h62 : _GEN_2730; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2732 = 8'hac == _t_T_18[31:24] ? 8'h91 : _GEN_2731; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2733 = 8'had == _t_T_18[31:24] ? 8'h95 : _GEN_2732; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2734 = 8'hae == _t_T_18[31:24] ? 8'he4 : _GEN_2733; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2735 = 8'haf == _t_T_18[31:24] ? 8'h79 : _GEN_2734; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2736 = 8'hb0 == _t_T_18[31:24] ? 8'he7 : _GEN_2735; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2737 = 8'hb1 == _t_T_18[31:24] ? 8'hc8 : _GEN_2736; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2738 = 8'hb2 == _t_T_18[31:24] ? 8'h37 : _GEN_2737; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2739 = 8'hb3 == _t_T_18[31:24] ? 8'h6d : _GEN_2738; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2740 = 8'hb4 == _t_T_18[31:24] ? 8'h8d : _GEN_2739; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2741 = 8'hb5 == _t_T_18[31:24] ? 8'hd5 : _GEN_2740; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2742 = 8'hb6 == _t_T_18[31:24] ? 8'h4e : _GEN_2741; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2743 = 8'hb7 == _t_T_18[31:24] ? 8'ha9 : _GEN_2742; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2744 = 8'hb8 == _t_T_18[31:24] ? 8'h6c : _GEN_2743; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2745 = 8'hb9 == _t_T_18[31:24] ? 8'h56 : _GEN_2744; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2746 = 8'hba == _t_T_18[31:24] ? 8'hf4 : _GEN_2745; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2747 = 8'hbb == _t_T_18[31:24] ? 8'hea : _GEN_2746; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2748 = 8'hbc == _t_T_18[31:24] ? 8'h65 : _GEN_2747; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2749 = 8'hbd == _t_T_18[31:24] ? 8'h7a : _GEN_2748; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2750 = 8'hbe == _t_T_18[31:24] ? 8'hae : _GEN_2749; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2751 = 8'hbf == _t_T_18[31:24] ? 8'h8 : _GEN_2750; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2752 = 8'hc0 == _t_T_18[31:24] ? 8'hba : _GEN_2751; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2753 = 8'hc1 == _t_T_18[31:24] ? 8'h78 : _GEN_2752; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2754 = 8'hc2 == _t_T_18[31:24] ? 8'h25 : _GEN_2753; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2755 = 8'hc3 == _t_T_18[31:24] ? 8'h2e : _GEN_2754; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2756 = 8'hc4 == _t_T_18[31:24] ? 8'h1c : _GEN_2755; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2757 = 8'hc5 == _t_T_18[31:24] ? 8'ha6 : _GEN_2756; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2758 = 8'hc6 == _t_T_18[31:24] ? 8'hb4 : _GEN_2757; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2759 = 8'hc7 == _t_T_18[31:24] ? 8'hc6 : _GEN_2758; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2760 = 8'hc8 == _t_T_18[31:24] ? 8'he8 : _GEN_2759; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2761 = 8'hc9 == _t_T_18[31:24] ? 8'hdd : _GEN_2760; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2762 = 8'hca == _t_T_18[31:24] ? 8'h74 : _GEN_2761; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2763 = 8'hcb == _t_T_18[31:24] ? 8'h1f : _GEN_2762; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2764 = 8'hcc == _t_T_18[31:24] ? 8'h4b : _GEN_2763; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2765 = 8'hcd == _t_T_18[31:24] ? 8'hbd : _GEN_2764; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2766 = 8'hce == _t_T_18[31:24] ? 8'h8b : _GEN_2765; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2767 = 8'hcf == _t_T_18[31:24] ? 8'h8a : _GEN_2766; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2768 = 8'hd0 == _t_T_18[31:24] ? 8'h70 : _GEN_2767; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2769 = 8'hd1 == _t_T_18[31:24] ? 8'h3e : _GEN_2768; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2770 = 8'hd2 == _t_T_18[31:24] ? 8'hb5 : _GEN_2769; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2771 = 8'hd3 == _t_T_18[31:24] ? 8'h66 : _GEN_2770; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2772 = 8'hd4 == _t_T_18[31:24] ? 8'h48 : _GEN_2771; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2773 = 8'hd5 == _t_T_18[31:24] ? 8'h3 : _GEN_2772; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2774 = 8'hd6 == _t_T_18[31:24] ? 8'hf6 : _GEN_2773; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2775 = 8'hd7 == _t_T_18[31:24] ? 8'he : _GEN_2774; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2776 = 8'hd8 == _t_T_18[31:24] ? 8'h61 : _GEN_2775; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2777 = 8'hd9 == _t_T_18[31:24] ? 8'h35 : _GEN_2776; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2778 = 8'hda == _t_T_18[31:24] ? 8'h57 : _GEN_2777; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2779 = 8'hdb == _t_T_18[31:24] ? 8'hb9 : _GEN_2778; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2780 = 8'hdc == _t_T_18[31:24] ? 8'h86 : _GEN_2779; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2781 = 8'hdd == _t_T_18[31:24] ? 8'hc1 : _GEN_2780; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2782 = 8'hde == _t_T_18[31:24] ? 8'h1d : _GEN_2781; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2783 = 8'hdf == _t_T_18[31:24] ? 8'h9e : _GEN_2782; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2784 = 8'he0 == _t_T_18[31:24] ? 8'he1 : _GEN_2783; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2785 = 8'he1 == _t_T_18[31:24] ? 8'hf8 : _GEN_2784; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2786 = 8'he2 == _t_T_18[31:24] ? 8'h98 : _GEN_2785; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2787 = 8'he3 == _t_T_18[31:24] ? 8'h11 : _GEN_2786; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2788 = 8'he4 == _t_T_18[31:24] ? 8'h69 : _GEN_2787; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2789 = 8'he5 == _t_T_18[31:24] ? 8'hd9 : _GEN_2788; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2790 = 8'he6 == _t_T_18[31:24] ? 8'h8e : _GEN_2789; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2791 = 8'he7 == _t_T_18[31:24] ? 8'h94 : _GEN_2790; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2792 = 8'he8 == _t_T_18[31:24] ? 8'h9b : _GEN_2791; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2793 = 8'he9 == _t_T_18[31:24] ? 8'h1e : _GEN_2792; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2794 = 8'hea == _t_T_18[31:24] ? 8'h87 : _GEN_2793; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2795 = 8'heb == _t_T_18[31:24] ? 8'he9 : _GEN_2794; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2796 = 8'hec == _t_T_18[31:24] ? 8'hce : _GEN_2795; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2797 = 8'hed == _t_T_18[31:24] ? 8'h55 : _GEN_2796; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2798 = 8'hee == _t_T_18[31:24] ? 8'h28 : _GEN_2797; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2799 = 8'hef == _t_T_18[31:24] ? 8'hdf : _GEN_2798; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2800 = 8'hf0 == _t_T_18[31:24] ? 8'h8c : _GEN_2799; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2801 = 8'hf1 == _t_T_18[31:24] ? 8'ha1 : _GEN_2800; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2802 = 8'hf2 == _t_T_18[31:24] ? 8'h89 : _GEN_2801; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2803 = 8'hf3 == _t_T_18[31:24] ? 8'hd : _GEN_2802; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2804 = 8'hf4 == _t_T_18[31:24] ? 8'hbf : _GEN_2803; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2805 = 8'hf5 == _t_T_18[31:24] ? 8'he6 : _GEN_2804; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2806 = 8'hf6 == _t_T_18[31:24] ? 8'h42 : _GEN_2805; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2807 = 8'hf7 == _t_T_18[31:24] ? 8'h68 : _GEN_2806; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2808 = 8'hf8 == _t_T_18[31:24] ? 8'h41 : _GEN_2807; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2809 = 8'hf9 == _t_T_18[31:24] ? 8'h99 : _GEN_2808; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2810 = 8'hfa == _t_T_18[31:24] ? 8'h2d : _GEN_2809; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2811 = 8'hfb == _t_T_18[31:24] ? 8'hf : _GEN_2810; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2812 = 8'hfc == _t_T_18[31:24] ? 8'hb0 : _GEN_2811; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2813 = 8'hfd == _t_T_18[31:24] ? 8'h54 : _GEN_2812; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2814 = 8'hfe == _t_T_18[31:24] ? 8'hbb : _GEN_2813; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2815 = 8'hff == _t_T_18[31:24] ? 8'h16 : _GEN_2814; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2817 = 8'h1 == _t_T_18[23:16] ? 8'h7c : 8'h63; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2818 = 8'h2 == _t_T_18[23:16] ? 8'h77 : _GEN_2817; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2819 = 8'h3 == _t_T_18[23:16] ? 8'h7b : _GEN_2818; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2820 = 8'h4 == _t_T_18[23:16] ? 8'hf2 : _GEN_2819; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2821 = 8'h5 == _t_T_18[23:16] ? 8'h6b : _GEN_2820; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2822 = 8'h6 == _t_T_18[23:16] ? 8'h6f : _GEN_2821; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2823 = 8'h7 == _t_T_18[23:16] ? 8'hc5 : _GEN_2822; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2824 = 8'h8 == _t_T_18[23:16] ? 8'h30 : _GEN_2823; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2825 = 8'h9 == _t_T_18[23:16] ? 8'h1 : _GEN_2824; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2826 = 8'ha == _t_T_18[23:16] ? 8'h67 : _GEN_2825; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2827 = 8'hb == _t_T_18[23:16] ? 8'h2b : _GEN_2826; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2828 = 8'hc == _t_T_18[23:16] ? 8'hfe : _GEN_2827; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2829 = 8'hd == _t_T_18[23:16] ? 8'hd7 : _GEN_2828; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2830 = 8'he == _t_T_18[23:16] ? 8'hab : _GEN_2829; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2831 = 8'hf == _t_T_18[23:16] ? 8'h76 : _GEN_2830; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2832 = 8'h10 == _t_T_18[23:16] ? 8'hca : _GEN_2831; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2833 = 8'h11 == _t_T_18[23:16] ? 8'h82 : _GEN_2832; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2834 = 8'h12 == _t_T_18[23:16] ? 8'hc9 : _GEN_2833; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2835 = 8'h13 == _t_T_18[23:16] ? 8'h7d : _GEN_2834; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2836 = 8'h14 == _t_T_18[23:16] ? 8'hfa : _GEN_2835; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2837 = 8'h15 == _t_T_18[23:16] ? 8'h59 : _GEN_2836; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2838 = 8'h16 == _t_T_18[23:16] ? 8'h47 : _GEN_2837; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2839 = 8'h17 == _t_T_18[23:16] ? 8'hf0 : _GEN_2838; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2840 = 8'h18 == _t_T_18[23:16] ? 8'had : _GEN_2839; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2841 = 8'h19 == _t_T_18[23:16] ? 8'hd4 : _GEN_2840; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2842 = 8'h1a == _t_T_18[23:16] ? 8'ha2 : _GEN_2841; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2843 = 8'h1b == _t_T_18[23:16] ? 8'haf : _GEN_2842; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2844 = 8'h1c == _t_T_18[23:16] ? 8'h9c : _GEN_2843; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2845 = 8'h1d == _t_T_18[23:16] ? 8'ha4 : _GEN_2844; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2846 = 8'h1e == _t_T_18[23:16] ? 8'h72 : _GEN_2845; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2847 = 8'h1f == _t_T_18[23:16] ? 8'hc0 : _GEN_2846; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2848 = 8'h20 == _t_T_18[23:16] ? 8'hb7 : _GEN_2847; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2849 = 8'h21 == _t_T_18[23:16] ? 8'hfd : _GEN_2848; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2850 = 8'h22 == _t_T_18[23:16] ? 8'h93 : _GEN_2849; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2851 = 8'h23 == _t_T_18[23:16] ? 8'h26 : _GEN_2850; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2852 = 8'h24 == _t_T_18[23:16] ? 8'h36 : _GEN_2851; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2853 = 8'h25 == _t_T_18[23:16] ? 8'h3f : _GEN_2852; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2854 = 8'h26 == _t_T_18[23:16] ? 8'hf7 : _GEN_2853; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2855 = 8'h27 == _t_T_18[23:16] ? 8'hcc : _GEN_2854; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2856 = 8'h28 == _t_T_18[23:16] ? 8'h34 : _GEN_2855; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2857 = 8'h29 == _t_T_18[23:16] ? 8'ha5 : _GEN_2856; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2858 = 8'h2a == _t_T_18[23:16] ? 8'he5 : _GEN_2857; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2859 = 8'h2b == _t_T_18[23:16] ? 8'hf1 : _GEN_2858; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2860 = 8'h2c == _t_T_18[23:16] ? 8'h71 : _GEN_2859; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2861 = 8'h2d == _t_T_18[23:16] ? 8'hd8 : _GEN_2860; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2862 = 8'h2e == _t_T_18[23:16] ? 8'h31 : _GEN_2861; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2863 = 8'h2f == _t_T_18[23:16] ? 8'h15 : _GEN_2862; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2864 = 8'h30 == _t_T_18[23:16] ? 8'h4 : _GEN_2863; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2865 = 8'h31 == _t_T_18[23:16] ? 8'hc7 : _GEN_2864; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2866 = 8'h32 == _t_T_18[23:16] ? 8'h23 : _GEN_2865; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2867 = 8'h33 == _t_T_18[23:16] ? 8'hc3 : _GEN_2866; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2868 = 8'h34 == _t_T_18[23:16] ? 8'h18 : _GEN_2867; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2869 = 8'h35 == _t_T_18[23:16] ? 8'h96 : _GEN_2868; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2870 = 8'h36 == _t_T_18[23:16] ? 8'h5 : _GEN_2869; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2871 = 8'h37 == _t_T_18[23:16] ? 8'h9a : _GEN_2870; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2872 = 8'h38 == _t_T_18[23:16] ? 8'h7 : _GEN_2871; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2873 = 8'h39 == _t_T_18[23:16] ? 8'h12 : _GEN_2872; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2874 = 8'h3a == _t_T_18[23:16] ? 8'h80 : _GEN_2873; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2875 = 8'h3b == _t_T_18[23:16] ? 8'he2 : _GEN_2874; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2876 = 8'h3c == _t_T_18[23:16] ? 8'heb : _GEN_2875; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2877 = 8'h3d == _t_T_18[23:16] ? 8'h27 : _GEN_2876; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2878 = 8'h3e == _t_T_18[23:16] ? 8'hb2 : _GEN_2877; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2879 = 8'h3f == _t_T_18[23:16] ? 8'h75 : _GEN_2878; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2880 = 8'h40 == _t_T_18[23:16] ? 8'h9 : _GEN_2879; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2881 = 8'h41 == _t_T_18[23:16] ? 8'h83 : _GEN_2880; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2882 = 8'h42 == _t_T_18[23:16] ? 8'h2c : _GEN_2881; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2883 = 8'h43 == _t_T_18[23:16] ? 8'h1a : _GEN_2882; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2884 = 8'h44 == _t_T_18[23:16] ? 8'h1b : _GEN_2883; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2885 = 8'h45 == _t_T_18[23:16] ? 8'h6e : _GEN_2884; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2886 = 8'h46 == _t_T_18[23:16] ? 8'h5a : _GEN_2885; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2887 = 8'h47 == _t_T_18[23:16] ? 8'ha0 : _GEN_2886; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2888 = 8'h48 == _t_T_18[23:16] ? 8'h52 : _GEN_2887; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2889 = 8'h49 == _t_T_18[23:16] ? 8'h3b : _GEN_2888; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2890 = 8'h4a == _t_T_18[23:16] ? 8'hd6 : _GEN_2889; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2891 = 8'h4b == _t_T_18[23:16] ? 8'hb3 : _GEN_2890; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2892 = 8'h4c == _t_T_18[23:16] ? 8'h29 : _GEN_2891; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2893 = 8'h4d == _t_T_18[23:16] ? 8'he3 : _GEN_2892; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2894 = 8'h4e == _t_T_18[23:16] ? 8'h2f : _GEN_2893; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2895 = 8'h4f == _t_T_18[23:16] ? 8'h84 : _GEN_2894; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2896 = 8'h50 == _t_T_18[23:16] ? 8'h53 : _GEN_2895; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2897 = 8'h51 == _t_T_18[23:16] ? 8'hd1 : _GEN_2896; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2898 = 8'h52 == _t_T_18[23:16] ? 8'h0 : _GEN_2897; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2899 = 8'h53 == _t_T_18[23:16] ? 8'hed : _GEN_2898; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2900 = 8'h54 == _t_T_18[23:16] ? 8'h20 : _GEN_2899; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2901 = 8'h55 == _t_T_18[23:16] ? 8'hfc : _GEN_2900; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2902 = 8'h56 == _t_T_18[23:16] ? 8'hb1 : _GEN_2901; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2903 = 8'h57 == _t_T_18[23:16] ? 8'h5b : _GEN_2902; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2904 = 8'h58 == _t_T_18[23:16] ? 8'h6a : _GEN_2903; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2905 = 8'h59 == _t_T_18[23:16] ? 8'hcb : _GEN_2904; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2906 = 8'h5a == _t_T_18[23:16] ? 8'hbe : _GEN_2905; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2907 = 8'h5b == _t_T_18[23:16] ? 8'h39 : _GEN_2906; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2908 = 8'h5c == _t_T_18[23:16] ? 8'h4a : _GEN_2907; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2909 = 8'h5d == _t_T_18[23:16] ? 8'h4c : _GEN_2908; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2910 = 8'h5e == _t_T_18[23:16] ? 8'h58 : _GEN_2909; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2911 = 8'h5f == _t_T_18[23:16] ? 8'hcf : _GEN_2910; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2912 = 8'h60 == _t_T_18[23:16] ? 8'hd0 : _GEN_2911; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2913 = 8'h61 == _t_T_18[23:16] ? 8'hef : _GEN_2912; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2914 = 8'h62 == _t_T_18[23:16] ? 8'haa : _GEN_2913; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2915 = 8'h63 == _t_T_18[23:16] ? 8'hfb : _GEN_2914; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2916 = 8'h64 == _t_T_18[23:16] ? 8'h43 : _GEN_2915; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2917 = 8'h65 == _t_T_18[23:16] ? 8'h4d : _GEN_2916; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2918 = 8'h66 == _t_T_18[23:16] ? 8'h33 : _GEN_2917; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2919 = 8'h67 == _t_T_18[23:16] ? 8'h85 : _GEN_2918; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2920 = 8'h68 == _t_T_18[23:16] ? 8'h45 : _GEN_2919; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2921 = 8'h69 == _t_T_18[23:16] ? 8'hf9 : _GEN_2920; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2922 = 8'h6a == _t_T_18[23:16] ? 8'h2 : _GEN_2921; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2923 = 8'h6b == _t_T_18[23:16] ? 8'h7f : _GEN_2922; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2924 = 8'h6c == _t_T_18[23:16] ? 8'h50 : _GEN_2923; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2925 = 8'h6d == _t_T_18[23:16] ? 8'h3c : _GEN_2924; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2926 = 8'h6e == _t_T_18[23:16] ? 8'h9f : _GEN_2925; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2927 = 8'h6f == _t_T_18[23:16] ? 8'ha8 : _GEN_2926; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2928 = 8'h70 == _t_T_18[23:16] ? 8'h51 : _GEN_2927; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2929 = 8'h71 == _t_T_18[23:16] ? 8'ha3 : _GEN_2928; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2930 = 8'h72 == _t_T_18[23:16] ? 8'h40 : _GEN_2929; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2931 = 8'h73 == _t_T_18[23:16] ? 8'h8f : _GEN_2930; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2932 = 8'h74 == _t_T_18[23:16] ? 8'h92 : _GEN_2931; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2933 = 8'h75 == _t_T_18[23:16] ? 8'h9d : _GEN_2932; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2934 = 8'h76 == _t_T_18[23:16] ? 8'h38 : _GEN_2933; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2935 = 8'h77 == _t_T_18[23:16] ? 8'hf5 : _GEN_2934; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2936 = 8'h78 == _t_T_18[23:16] ? 8'hbc : _GEN_2935; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2937 = 8'h79 == _t_T_18[23:16] ? 8'hb6 : _GEN_2936; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2938 = 8'h7a == _t_T_18[23:16] ? 8'hda : _GEN_2937; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2939 = 8'h7b == _t_T_18[23:16] ? 8'h21 : _GEN_2938; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2940 = 8'h7c == _t_T_18[23:16] ? 8'h10 : _GEN_2939; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2941 = 8'h7d == _t_T_18[23:16] ? 8'hff : _GEN_2940; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2942 = 8'h7e == _t_T_18[23:16] ? 8'hf3 : _GEN_2941; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2943 = 8'h7f == _t_T_18[23:16] ? 8'hd2 : _GEN_2942; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2944 = 8'h80 == _t_T_18[23:16] ? 8'hcd : _GEN_2943; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2945 = 8'h81 == _t_T_18[23:16] ? 8'hc : _GEN_2944; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2946 = 8'h82 == _t_T_18[23:16] ? 8'h13 : _GEN_2945; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2947 = 8'h83 == _t_T_18[23:16] ? 8'hec : _GEN_2946; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2948 = 8'h84 == _t_T_18[23:16] ? 8'h5f : _GEN_2947; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2949 = 8'h85 == _t_T_18[23:16] ? 8'h97 : _GEN_2948; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2950 = 8'h86 == _t_T_18[23:16] ? 8'h44 : _GEN_2949; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2951 = 8'h87 == _t_T_18[23:16] ? 8'h17 : _GEN_2950; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2952 = 8'h88 == _t_T_18[23:16] ? 8'hc4 : _GEN_2951; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2953 = 8'h89 == _t_T_18[23:16] ? 8'ha7 : _GEN_2952; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2954 = 8'h8a == _t_T_18[23:16] ? 8'h7e : _GEN_2953; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2955 = 8'h8b == _t_T_18[23:16] ? 8'h3d : _GEN_2954; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2956 = 8'h8c == _t_T_18[23:16] ? 8'h64 : _GEN_2955; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2957 = 8'h8d == _t_T_18[23:16] ? 8'h5d : _GEN_2956; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2958 = 8'h8e == _t_T_18[23:16] ? 8'h19 : _GEN_2957; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2959 = 8'h8f == _t_T_18[23:16] ? 8'h73 : _GEN_2958; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2960 = 8'h90 == _t_T_18[23:16] ? 8'h60 : _GEN_2959; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2961 = 8'h91 == _t_T_18[23:16] ? 8'h81 : _GEN_2960; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2962 = 8'h92 == _t_T_18[23:16] ? 8'h4f : _GEN_2961; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2963 = 8'h93 == _t_T_18[23:16] ? 8'hdc : _GEN_2962; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2964 = 8'h94 == _t_T_18[23:16] ? 8'h22 : _GEN_2963; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2965 = 8'h95 == _t_T_18[23:16] ? 8'h2a : _GEN_2964; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2966 = 8'h96 == _t_T_18[23:16] ? 8'h90 : _GEN_2965; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2967 = 8'h97 == _t_T_18[23:16] ? 8'h88 : _GEN_2966; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2968 = 8'h98 == _t_T_18[23:16] ? 8'h46 : _GEN_2967; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2969 = 8'h99 == _t_T_18[23:16] ? 8'hee : _GEN_2968; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2970 = 8'h9a == _t_T_18[23:16] ? 8'hb8 : _GEN_2969; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2971 = 8'h9b == _t_T_18[23:16] ? 8'h14 : _GEN_2970; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2972 = 8'h9c == _t_T_18[23:16] ? 8'hde : _GEN_2971; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2973 = 8'h9d == _t_T_18[23:16] ? 8'h5e : _GEN_2972; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2974 = 8'h9e == _t_T_18[23:16] ? 8'hb : _GEN_2973; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2975 = 8'h9f == _t_T_18[23:16] ? 8'hdb : _GEN_2974; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2976 = 8'ha0 == _t_T_18[23:16] ? 8'he0 : _GEN_2975; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2977 = 8'ha1 == _t_T_18[23:16] ? 8'h32 : _GEN_2976; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2978 = 8'ha2 == _t_T_18[23:16] ? 8'h3a : _GEN_2977; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2979 = 8'ha3 == _t_T_18[23:16] ? 8'ha : _GEN_2978; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2980 = 8'ha4 == _t_T_18[23:16] ? 8'h49 : _GEN_2979; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2981 = 8'ha5 == _t_T_18[23:16] ? 8'h6 : _GEN_2980; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2982 = 8'ha6 == _t_T_18[23:16] ? 8'h24 : _GEN_2981; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2983 = 8'ha7 == _t_T_18[23:16] ? 8'h5c : _GEN_2982; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2984 = 8'ha8 == _t_T_18[23:16] ? 8'hc2 : _GEN_2983; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2985 = 8'ha9 == _t_T_18[23:16] ? 8'hd3 : _GEN_2984; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2986 = 8'haa == _t_T_18[23:16] ? 8'hac : _GEN_2985; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2987 = 8'hab == _t_T_18[23:16] ? 8'h62 : _GEN_2986; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2988 = 8'hac == _t_T_18[23:16] ? 8'h91 : _GEN_2987; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2989 = 8'had == _t_T_18[23:16] ? 8'h95 : _GEN_2988; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2990 = 8'hae == _t_T_18[23:16] ? 8'he4 : _GEN_2989; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2991 = 8'haf == _t_T_18[23:16] ? 8'h79 : _GEN_2990; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2992 = 8'hb0 == _t_T_18[23:16] ? 8'he7 : _GEN_2991; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2993 = 8'hb1 == _t_T_18[23:16] ? 8'hc8 : _GEN_2992; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2994 = 8'hb2 == _t_T_18[23:16] ? 8'h37 : _GEN_2993; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2995 = 8'hb3 == _t_T_18[23:16] ? 8'h6d : _GEN_2994; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2996 = 8'hb4 == _t_T_18[23:16] ? 8'h8d : _GEN_2995; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2997 = 8'hb5 == _t_T_18[23:16] ? 8'hd5 : _GEN_2996; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2998 = 8'hb6 == _t_T_18[23:16] ? 8'h4e : _GEN_2997; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_2999 = 8'hb7 == _t_T_18[23:16] ? 8'ha9 : _GEN_2998; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3000 = 8'hb8 == _t_T_18[23:16] ? 8'h6c : _GEN_2999; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3001 = 8'hb9 == _t_T_18[23:16] ? 8'h56 : _GEN_3000; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3002 = 8'hba == _t_T_18[23:16] ? 8'hf4 : _GEN_3001; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3003 = 8'hbb == _t_T_18[23:16] ? 8'hea : _GEN_3002; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3004 = 8'hbc == _t_T_18[23:16] ? 8'h65 : _GEN_3003; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3005 = 8'hbd == _t_T_18[23:16] ? 8'h7a : _GEN_3004; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3006 = 8'hbe == _t_T_18[23:16] ? 8'hae : _GEN_3005; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3007 = 8'hbf == _t_T_18[23:16] ? 8'h8 : _GEN_3006; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3008 = 8'hc0 == _t_T_18[23:16] ? 8'hba : _GEN_3007; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3009 = 8'hc1 == _t_T_18[23:16] ? 8'h78 : _GEN_3008; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3010 = 8'hc2 == _t_T_18[23:16] ? 8'h25 : _GEN_3009; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3011 = 8'hc3 == _t_T_18[23:16] ? 8'h2e : _GEN_3010; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3012 = 8'hc4 == _t_T_18[23:16] ? 8'h1c : _GEN_3011; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3013 = 8'hc5 == _t_T_18[23:16] ? 8'ha6 : _GEN_3012; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3014 = 8'hc6 == _t_T_18[23:16] ? 8'hb4 : _GEN_3013; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3015 = 8'hc7 == _t_T_18[23:16] ? 8'hc6 : _GEN_3014; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3016 = 8'hc8 == _t_T_18[23:16] ? 8'he8 : _GEN_3015; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3017 = 8'hc9 == _t_T_18[23:16] ? 8'hdd : _GEN_3016; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3018 = 8'hca == _t_T_18[23:16] ? 8'h74 : _GEN_3017; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3019 = 8'hcb == _t_T_18[23:16] ? 8'h1f : _GEN_3018; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3020 = 8'hcc == _t_T_18[23:16] ? 8'h4b : _GEN_3019; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3021 = 8'hcd == _t_T_18[23:16] ? 8'hbd : _GEN_3020; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3022 = 8'hce == _t_T_18[23:16] ? 8'h8b : _GEN_3021; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3023 = 8'hcf == _t_T_18[23:16] ? 8'h8a : _GEN_3022; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3024 = 8'hd0 == _t_T_18[23:16] ? 8'h70 : _GEN_3023; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3025 = 8'hd1 == _t_T_18[23:16] ? 8'h3e : _GEN_3024; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3026 = 8'hd2 == _t_T_18[23:16] ? 8'hb5 : _GEN_3025; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3027 = 8'hd3 == _t_T_18[23:16] ? 8'h66 : _GEN_3026; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3028 = 8'hd4 == _t_T_18[23:16] ? 8'h48 : _GEN_3027; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3029 = 8'hd5 == _t_T_18[23:16] ? 8'h3 : _GEN_3028; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3030 = 8'hd6 == _t_T_18[23:16] ? 8'hf6 : _GEN_3029; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3031 = 8'hd7 == _t_T_18[23:16] ? 8'he : _GEN_3030; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3032 = 8'hd8 == _t_T_18[23:16] ? 8'h61 : _GEN_3031; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3033 = 8'hd9 == _t_T_18[23:16] ? 8'h35 : _GEN_3032; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3034 = 8'hda == _t_T_18[23:16] ? 8'h57 : _GEN_3033; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3035 = 8'hdb == _t_T_18[23:16] ? 8'hb9 : _GEN_3034; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3036 = 8'hdc == _t_T_18[23:16] ? 8'h86 : _GEN_3035; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3037 = 8'hdd == _t_T_18[23:16] ? 8'hc1 : _GEN_3036; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3038 = 8'hde == _t_T_18[23:16] ? 8'h1d : _GEN_3037; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3039 = 8'hdf == _t_T_18[23:16] ? 8'h9e : _GEN_3038; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3040 = 8'he0 == _t_T_18[23:16] ? 8'he1 : _GEN_3039; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3041 = 8'he1 == _t_T_18[23:16] ? 8'hf8 : _GEN_3040; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3042 = 8'he2 == _t_T_18[23:16] ? 8'h98 : _GEN_3041; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3043 = 8'he3 == _t_T_18[23:16] ? 8'h11 : _GEN_3042; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3044 = 8'he4 == _t_T_18[23:16] ? 8'h69 : _GEN_3043; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3045 = 8'he5 == _t_T_18[23:16] ? 8'hd9 : _GEN_3044; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3046 = 8'he6 == _t_T_18[23:16] ? 8'h8e : _GEN_3045; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3047 = 8'he7 == _t_T_18[23:16] ? 8'h94 : _GEN_3046; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3048 = 8'he8 == _t_T_18[23:16] ? 8'h9b : _GEN_3047; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3049 = 8'he9 == _t_T_18[23:16] ? 8'h1e : _GEN_3048; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3050 = 8'hea == _t_T_18[23:16] ? 8'h87 : _GEN_3049; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3051 = 8'heb == _t_T_18[23:16] ? 8'he9 : _GEN_3050; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3052 = 8'hec == _t_T_18[23:16] ? 8'hce : _GEN_3051; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3053 = 8'hed == _t_T_18[23:16] ? 8'h55 : _GEN_3052; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3054 = 8'hee == _t_T_18[23:16] ? 8'h28 : _GEN_3053; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3055 = 8'hef == _t_T_18[23:16] ? 8'hdf : _GEN_3054; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3056 = 8'hf0 == _t_T_18[23:16] ? 8'h8c : _GEN_3055; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3057 = 8'hf1 == _t_T_18[23:16] ? 8'ha1 : _GEN_3056; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3058 = 8'hf2 == _t_T_18[23:16] ? 8'h89 : _GEN_3057; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3059 = 8'hf3 == _t_T_18[23:16] ? 8'hd : _GEN_3058; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3060 = 8'hf4 == _t_T_18[23:16] ? 8'hbf : _GEN_3059; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3061 = 8'hf5 == _t_T_18[23:16] ? 8'he6 : _GEN_3060; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3062 = 8'hf6 == _t_T_18[23:16] ? 8'h42 : _GEN_3061; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3063 = 8'hf7 == _t_T_18[23:16] ? 8'h68 : _GEN_3062; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3064 = 8'hf8 == _t_T_18[23:16] ? 8'h41 : _GEN_3063; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3065 = 8'hf9 == _t_T_18[23:16] ? 8'h99 : _GEN_3064; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3066 = 8'hfa == _t_T_18[23:16] ? 8'h2d : _GEN_3065; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3067 = 8'hfb == _t_T_18[23:16] ? 8'hf : _GEN_3066; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3068 = 8'hfc == _t_T_18[23:16] ? 8'hb0 : _GEN_3067; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3069 = 8'hfd == _t_T_18[23:16] ? 8'h54 : _GEN_3068; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3070 = 8'hfe == _t_T_18[23:16] ? 8'hbb : _GEN_3069; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3071 = 8'hff == _t_T_18[23:16] ? 8'h16 : _GEN_3070; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [31:0] _t_T_23 = {_GEN_2815,_GEN_3071,_GEN_2303,_GEN_2559}; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:8]
  wire [31:0] t_2 = _t_T_23 ^ 32'h4000000; // @[src/main/scala/crypto/aes/KeySchedule.scala 59:32]
  wire [31:0] w_12 = w_8 ^ t_2; // @[src/main/scala/crypto/aes/KeySchedule.scala 63:21]
  wire [31:0] w_13 = w_9 ^ w_12; // @[src/main/scala/crypto/aes/KeySchedule.scala 63:21]
  wire [31:0] w_14 = w_10 ^ w_13; // @[src/main/scala/crypto/aes/KeySchedule.scala 63:21]
  wire [31:0] w_15 = w_11 ^ w_14; // @[src/main/scala/crypto/aes/KeySchedule.scala 63:21]
  wire [31:0] _t_T_26 = {w_15[23:0],w_15[31:24]}; // @[src/main/scala/crypto/aes/KeySchedule.scala 23:43]
  wire [7:0] _GEN_3073 = 8'h1 == _t_T_26[15:8] ? 8'h7c : 8'h63; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3074 = 8'h2 == _t_T_26[15:8] ? 8'h77 : _GEN_3073; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3075 = 8'h3 == _t_T_26[15:8] ? 8'h7b : _GEN_3074; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3076 = 8'h4 == _t_T_26[15:8] ? 8'hf2 : _GEN_3075; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3077 = 8'h5 == _t_T_26[15:8] ? 8'h6b : _GEN_3076; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3078 = 8'h6 == _t_T_26[15:8] ? 8'h6f : _GEN_3077; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3079 = 8'h7 == _t_T_26[15:8] ? 8'hc5 : _GEN_3078; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3080 = 8'h8 == _t_T_26[15:8] ? 8'h30 : _GEN_3079; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3081 = 8'h9 == _t_T_26[15:8] ? 8'h1 : _GEN_3080; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3082 = 8'ha == _t_T_26[15:8] ? 8'h67 : _GEN_3081; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3083 = 8'hb == _t_T_26[15:8] ? 8'h2b : _GEN_3082; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3084 = 8'hc == _t_T_26[15:8] ? 8'hfe : _GEN_3083; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3085 = 8'hd == _t_T_26[15:8] ? 8'hd7 : _GEN_3084; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3086 = 8'he == _t_T_26[15:8] ? 8'hab : _GEN_3085; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3087 = 8'hf == _t_T_26[15:8] ? 8'h76 : _GEN_3086; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3088 = 8'h10 == _t_T_26[15:8] ? 8'hca : _GEN_3087; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3089 = 8'h11 == _t_T_26[15:8] ? 8'h82 : _GEN_3088; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3090 = 8'h12 == _t_T_26[15:8] ? 8'hc9 : _GEN_3089; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3091 = 8'h13 == _t_T_26[15:8] ? 8'h7d : _GEN_3090; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3092 = 8'h14 == _t_T_26[15:8] ? 8'hfa : _GEN_3091; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3093 = 8'h15 == _t_T_26[15:8] ? 8'h59 : _GEN_3092; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3094 = 8'h16 == _t_T_26[15:8] ? 8'h47 : _GEN_3093; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3095 = 8'h17 == _t_T_26[15:8] ? 8'hf0 : _GEN_3094; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3096 = 8'h18 == _t_T_26[15:8] ? 8'had : _GEN_3095; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3097 = 8'h19 == _t_T_26[15:8] ? 8'hd4 : _GEN_3096; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3098 = 8'h1a == _t_T_26[15:8] ? 8'ha2 : _GEN_3097; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3099 = 8'h1b == _t_T_26[15:8] ? 8'haf : _GEN_3098; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3100 = 8'h1c == _t_T_26[15:8] ? 8'h9c : _GEN_3099; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3101 = 8'h1d == _t_T_26[15:8] ? 8'ha4 : _GEN_3100; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3102 = 8'h1e == _t_T_26[15:8] ? 8'h72 : _GEN_3101; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3103 = 8'h1f == _t_T_26[15:8] ? 8'hc0 : _GEN_3102; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3104 = 8'h20 == _t_T_26[15:8] ? 8'hb7 : _GEN_3103; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3105 = 8'h21 == _t_T_26[15:8] ? 8'hfd : _GEN_3104; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3106 = 8'h22 == _t_T_26[15:8] ? 8'h93 : _GEN_3105; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3107 = 8'h23 == _t_T_26[15:8] ? 8'h26 : _GEN_3106; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3108 = 8'h24 == _t_T_26[15:8] ? 8'h36 : _GEN_3107; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3109 = 8'h25 == _t_T_26[15:8] ? 8'h3f : _GEN_3108; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3110 = 8'h26 == _t_T_26[15:8] ? 8'hf7 : _GEN_3109; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3111 = 8'h27 == _t_T_26[15:8] ? 8'hcc : _GEN_3110; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3112 = 8'h28 == _t_T_26[15:8] ? 8'h34 : _GEN_3111; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3113 = 8'h29 == _t_T_26[15:8] ? 8'ha5 : _GEN_3112; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3114 = 8'h2a == _t_T_26[15:8] ? 8'he5 : _GEN_3113; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3115 = 8'h2b == _t_T_26[15:8] ? 8'hf1 : _GEN_3114; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3116 = 8'h2c == _t_T_26[15:8] ? 8'h71 : _GEN_3115; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3117 = 8'h2d == _t_T_26[15:8] ? 8'hd8 : _GEN_3116; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3118 = 8'h2e == _t_T_26[15:8] ? 8'h31 : _GEN_3117; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3119 = 8'h2f == _t_T_26[15:8] ? 8'h15 : _GEN_3118; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3120 = 8'h30 == _t_T_26[15:8] ? 8'h4 : _GEN_3119; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3121 = 8'h31 == _t_T_26[15:8] ? 8'hc7 : _GEN_3120; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3122 = 8'h32 == _t_T_26[15:8] ? 8'h23 : _GEN_3121; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3123 = 8'h33 == _t_T_26[15:8] ? 8'hc3 : _GEN_3122; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3124 = 8'h34 == _t_T_26[15:8] ? 8'h18 : _GEN_3123; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3125 = 8'h35 == _t_T_26[15:8] ? 8'h96 : _GEN_3124; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3126 = 8'h36 == _t_T_26[15:8] ? 8'h5 : _GEN_3125; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3127 = 8'h37 == _t_T_26[15:8] ? 8'h9a : _GEN_3126; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3128 = 8'h38 == _t_T_26[15:8] ? 8'h7 : _GEN_3127; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3129 = 8'h39 == _t_T_26[15:8] ? 8'h12 : _GEN_3128; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3130 = 8'h3a == _t_T_26[15:8] ? 8'h80 : _GEN_3129; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3131 = 8'h3b == _t_T_26[15:8] ? 8'he2 : _GEN_3130; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3132 = 8'h3c == _t_T_26[15:8] ? 8'heb : _GEN_3131; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3133 = 8'h3d == _t_T_26[15:8] ? 8'h27 : _GEN_3132; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3134 = 8'h3e == _t_T_26[15:8] ? 8'hb2 : _GEN_3133; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3135 = 8'h3f == _t_T_26[15:8] ? 8'h75 : _GEN_3134; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3136 = 8'h40 == _t_T_26[15:8] ? 8'h9 : _GEN_3135; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3137 = 8'h41 == _t_T_26[15:8] ? 8'h83 : _GEN_3136; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3138 = 8'h42 == _t_T_26[15:8] ? 8'h2c : _GEN_3137; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3139 = 8'h43 == _t_T_26[15:8] ? 8'h1a : _GEN_3138; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3140 = 8'h44 == _t_T_26[15:8] ? 8'h1b : _GEN_3139; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3141 = 8'h45 == _t_T_26[15:8] ? 8'h6e : _GEN_3140; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3142 = 8'h46 == _t_T_26[15:8] ? 8'h5a : _GEN_3141; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3143 = 8'h47 == _t_T_26[15:8] ? 8'ha0 : _GEN_3142; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3144 = 8'h48 == _t_T_26[15:8] ? 8'h52 : _GEN_3143; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3145 = 8'h49 == _t_T_26[15:8] ? 8'h3b : _GEN_3144; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3146 = 8'h4a == _t_T_26[15:8] ? 8'hd6 : _GEN_3145; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3147 = 8'h4b == _t_T_26[15:8] ? 8'hb3 : _GEN_3146; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3148 = 8'h4c == _t_T_26[15:8] ? 8'h29 : _GEN_3147; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3149 = 8'h4d == _t_T_26[15:8] ? 8'he3 : _GEN_3148; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3150 = 8'h4e == _t_T_26[15:8] ? 8'h2f : _GEN_3149; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3151 = 8'h4f == _t_T_26[15:8] ? 8'h84 : _GEN_3150; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3152 = 8'h50 == _t_T_26[15:8] ? 8'h53 : _GEN_3151; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3153 = 8'h51 == _t_T_26[15:8] ? 8'hd1 : _GEN_3152; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3154 = 8'h52 == _t_T_26[15:8] ? 8'h0 : _GEN_3153; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3155 = 8'h53 == _t_T_26[15:8] ? 8'hed : _GEN_3154; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3156 = 8'h54 == _t_T_26[15:8] ? 8'h20 : _GEN_3155; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3157 = 8'h55 == _t_T_26[15:8] ? 8'hfc : _GEN_3156; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3158 = 8'h56 == _t_T_26[15:8] ? 8'hb1 : _GEN_3157; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3159 = 8'h57 == _t_T_26[15:8] ? 8'h5b : _GEN_3158; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3160 = 8'h58 == _t_T_26[15:8] ? 8'h6a : _GEN_3159; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3161 = 8'h59 == _t_T_26[15:8] ? 8'hcb : _GEN_3160; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3162 = 8'h5a == _t_T_26[15:8] ? 8'hbe : _GEN_3161; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3163 = 8'h5b == _t_T_26[15:8] ? 8'h39 : _GEN_3162; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3164 = 8'h5c == _t_T_26[15:8] ? 8'h4a : _GEN_3163; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3165 = 8'h5d == _t_T_26[15:8] ? 8'h4c : _GEN_3164; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3166 = 8'h5e == _t_T_26[15:8] ? 8'h58 : _GEN_3165; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3167 = 8'h5f == _t_T_26[15:8] ? 8'hcf : _GEN_3166; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3168 = 8'h60 == _t_T_26[15:8] ? 8'hd0 : _GEN_3167; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3169 = 8'h61 == _t_T_26[15:8] ? 8'hef : _GEN_3168; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3170 = 8'h62 == _t_T_26[15:8] ? 8'haa : _GEN_3169; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3171 = 8'h63 == _t_T_26[15:8] ? 8'hfb : _GEN_3170; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3172 = 8'h64 == _t_T_26[15:8] ? 8'h43 : _GEN_3171; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3173 = 8'h65 == _t_T_26[15:8] ? 8'h4d : _GEN_3172; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3174 = 8'h66 == _t_T_26[15:8] ? 8'h33 : _GEN_3173; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3175 = 8'h67 == _t_T_26[15:8] ? 8'h85 : _GEN_3174; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3176 = 8'h68 == _t_T_26[15:8] ? 8'h45 : _GEN_3175; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3177 = 8'h69 == _t_T_26[15:8] ? 8'hf9 : _GEN_3176; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3178 = 8'h6a == _t_T_26[15:8] ? 8'h2 : _GEN_3177; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3179 = 8'h6b == _t_T_26[15:8] ? 8'h7f : _GEN_3178; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3180 = 8'h6c == _t_T_26[15:8] ? 8'h50 : _GEN_3179; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3181 = 8'h6d == _t_T_26[15:8] ? 8'h3c : _GEN_3180; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3182 = 8'h6e == _t_T_26[15:8] ? 8'h9f : _GEN_3181; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3183 = 8'h6f == _t_T_26[15:8] ? 8'ha8 : _GEN_3182; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3184 = 8'h70 == _t_T_26[15:8] ? 8'h51 : _GEN_3183; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3185 = 8'h71 == _t_T_26[15:8] ? 8'ha3 : _GEN_3184; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3186 = 8'h72 == _t_T_26[15:8] ? 8'h40 : _GEN_3185; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3187 = 8'h73 == _t_T_26[15:8] ? 8'h8f : _GEN_3186; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3188 = 8'h74 == _t_T_26[15:8] ? 8'h92 : _GEN_3187; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3189 = 8'h75 == _t_T_26[15:8] ? 8'h9d : _GEN_3188; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3190 = 8'h76 == _t_T_26[15:8] ? 8'h38 : _GEN_3189; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3191 = 8'h77 == _t_T_26[15:8] ? 8'hf5 : _GEN_3190; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3192 = 8'h78 == _t_T_26[15:8] ? 8'hbc : _GEN_3191; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3193 = 8'h79 == _t_T_26[15:8] ? 8'hb6 : _GEN_3192; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3194 = 8'h7a == _t_T_26[15:8] ? 8'hda : _GEN_3193; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3195 = 8'h7b == _t_T_26[15:8] ? 8'h21 : _GEN_3194; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3196 = 8'h7c == _t_T_26[15:8] ? 8'h10 : _GEN_3195; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3197 = 8'h7d == _t_T_26[15:8] ? 8'hff : _GEN_3196; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3198 = 8'h7e == _t_T_26[15:8] ? 8'hf3 : _GEN_3197; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3199 = 8'h7f == _t_T_26[15:8] ? 8'hd2 : _GEN_3198; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3200 = 8'h80 == _t_T_26[15:8] ? 8'hcd : _GEN_3199; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3201 = 8'h81 == _t_T_26[15:8] ? 8'hc : _GEN_3200; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3202 = 8'h82 == _t_T_26[15:8] ? 8'h13 : _GEN_3201; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3203 = 8'h83 == _t_T_26[15:8] ? 8'hec : _GEN_3202; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3204 = 8'h84 == _t_T_26[15:8] ? 8'h5f : _GEN_3203; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3205 = 8'h85 == _t_T_26[15:8] ? 8'h97 : _GEN_3204; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3206 = 8'h86 == _t_T_26[15:8] ? 8'h44 : _GEN_3205; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3207 = 8'h87 == _t_T_26[15:8] ? 8'h17 : _GEN_3206; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3208 = 8'h88 == _t_T_26[15:8] ? 8'hc4 : _GEN_3207; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3209 = 8'h89 == _t_T_26[15:8] ? 8'ha7 : _GEN_3208; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3210 = 8'h8a == _t_T_26[15:8] ? 8'h7e : _GEN_3209; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3211 = 8'h8b == _t_T_26[15:8] ? 8'h3d : _GEN_3210; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3212 = 8'h8c == _t_T_26[15:8] ? 8'h64 : _GEN_3211; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3213 = 8'h8d == _t_T_26[15:8] ? 8'h5d : _GEN_3212; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3214 = 8'h8e == _t_T_26[15:8] ? 8'h19 : _GEN_3213; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3215 = 8'h8f == _t_T_26[15:8] ? 8'h73 : _GEN_3214; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3216 = 8'h90 == _t_T_26[15:8] ? 8'h60 : _GEN_3215; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3217 = 8'h91 == _t_T_26[15:8] ? 8'h81 : _GEN_3216; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3218 = 8'h92 == _t_T_26[15:8] ? 8'h4f : _GEN_3217; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3219 = 8'h93 == _t_T_26[15:8] ? 8'hdc : _GEN_3218; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3220 = 8'h94 == _t_T_26[15:8] ? 8'h22 : _GEN_3219; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3221 = 8'h95 == _t_T_26[15:8] ? 8'h2a : _GEN_3220; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3222 = 8'h96 == _t_T_26[15:8] ? 8'h90 : _GEN_3221; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3223 = 8'h97 == _t_T_26[15:8] ? 8'h88 : _GEN_3222; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3224 = 8'h98 == _t_T_26[15:8] ? 8'h46 : _GEN_3223; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3225 = 8'h99 == _t_T_26[15:8] ? 8'hee : _GEN_3224; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3226 = 8'h9a == _t_T_26[15:8] ? 8'hb8 : _GEN_3225; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3227 = 8'h9b == _t_T_26[15:8] ? 8'h14 : _GEN_3226; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3228 = 8'h9c == _t_T_26[15:8] ? 8'hde : _GEN_3227; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3229 = 8'h9d == _t_T_26[15:8] ? 8'h5e : _GEN_3228; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3230 = 8'h9e == _t_T_26[15:8] ? 8'hb : _GEN_3229; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3231 = 8'h9f == _t_T_26[15:8] ? 8'hdb : _GEN_3230; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3232 = 8'ha0 == _t_T_26[15:8] ? 8'he0 : _GEN_3231; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3233 = 8'ha1 == _t_T_26[15:8] ? 8'h32 : _GEN_3232; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3234 = 8'ha2 == _t_T_26[15:8] ? 8'h3a : _GEN_3233; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3235 = 8'ha3 == _t_T_26[15:8] ? 8'ha : _GEN_3234; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3236 = 8'ha4 == _t_T_26[15:8] ? 8'h49 : _GEN_3235; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3237 = 8'ha5 == _t_T_26[15:8] ? 8'h6 : _GEN_3236; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3238 = 8'ha6 == _t_T_26[15:8] ? 8'h24 : _GEN_3237; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3239 = 8'ha7 == _t_T_26[15:8] ? 8'h5c : _GEN_3238; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3240 = 8'ha8 == _t_T_26[15:8] ? 8'hc2 : _GEN_3239; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3241 = 8'ha9 == _t_T_26[15:8] ? 8'hd3 : _GEN_3240; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3242 = 8'haa == _t_T_26[15:8] ? 8'hac : _GEN_3241; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3243 = 8'hab == _t_T_26[15:8] ? 8'h62 : _GEN_3242; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3244 = 8'hac == _t_T_26[15:8] ? 8'h91 : _GEN_3243; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3245 = 8'had == _t_T_26[15:8] ? 8'h95 : _GEN_3244; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3246 = 8'hae == _t_T_26[15:8] ? 8'he4 : _GEN_3245; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3247 = 8'haf == _t_T_26[15:8] ? 8'h79 : _GEN_3246; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3248 = 8'hb0 == _t_T_26[15:8] ? 8'he7 : _GEN_3247; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3249 = 8'hb1 == _t_T_26[15:8] ? 8'hc8 : _GEN_3248; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3250 = 8'hb2 == _t_T_26[15:8] ? 8'h37 : _GEN_3249; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3251 = 8'hb3 == _t_T_26[15:8] ? 8'h6d : _GEN_3250; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3252 = 8'hb4 == _t_T_26[15:8] ? 8'h8d : _GEN_3251; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3253 = 8'hb5 == _t_T_26[15:8] ? 8'hd5 : _GEN_3252; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3254 = 8'hb6 == _t_T_26[15:8] ? 8'h4e : _GEN_3253; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3255 = 8'hb7 == _t_T_26[15:8] ? 8'ha9 : _GEN_3254; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3256 = 8'hb8 == _t_T_26[15:8] ? 8'h6c : _GEN_3255; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3257 = 8'hb9 == _t_T_26[15:8] ? 8'h56 : _GEN_3256; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3258 = 8'hba == _t_T_26[15:8] ? 8'hf4 : _GEN_3257; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3259 = 8'hbb == _t_T_26[15:8] ? 8'hea : _GEN_3258; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3260 = 8'hbc == _t_T_26[15:8] ? 8'h65 : _GEN_3259; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3261 = 8'hbd == _t_T_26[15:8] ? 8'h7a : _GEN_3260; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3262 = 8'hbe == _t_T_26[15:8] ? 8'hae : _GEN_3261; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3263 = 8'hbf == _t_T_26[15:8] ? 8'h8 : _GEN_3262; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3264 = 8'hc0 == _t_T_26[15:8] ? 8'hba : _GEN_3263; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3265 = 8'hc1 == _t_T_26[15:8] ? 8'h78 : _GEN_3264; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3266 = 8'hc2 == _t_T_26[15:8] ? 8'h25 : _GEN_3265; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3267 = 8'hc3 == _t_T_26[15:8] ? 8'h2e : _GEN_3266; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3268 = 8'hc4 == _t_T_26[15:8] ? 8'h1c : _GEN_3267; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3269 = 8'hc5 == _t_T_26[15:8] ? 8'ha6 : _GEN_3268; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3270 = 8'hc6 == _t_T_26[15:8] ? 8'hb4 : _GEN_3269; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3271 = 8'hc7 == _t_T_26[15:8] ? 8'hc6 : _GEN_3270; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3272 = 8'hc8 == _t_T_26[15:8] ? 8'he8 : _GEN_3271; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3273 = 8'hc9 == _t_T_26[15:8] ? 8'hdd : _GEN_3272; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3274 = 8'hca == _t_T_26[15:8] ? 8'h74 : _GEN_3273; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3275 = 8'hcb == _t_T_26[15:8] ? 8'h1f : _GEN_3274; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3276 = 8'hcc == _t_T_26[15:8] ? 8'h4b : _GEN_3275; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3277 = 8'hcd == _t_T_26[15:8] ? 8'hbd : _GEN_3276; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3278 = 8'hce == _t_T_26[15:8] ? 8'h8b : _GEN_3277; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3279 = 8'hcf == _t_T_26[15:8] ? 8'h8a : _GEN_3278; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3280 = 8'hd0 == _t_T_26[15:8] ? 8'h70 : _GEN_3279; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3281 = 8'hd1 == _t_T_26[15:8] ? 8'h3e : _GEN_3280; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3282 = 8'hd2 == _t_T_26[15:8] ? 8'hb5 : _GEN_3281; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3283 = 8'hd3 == _t_T_26[15:8] ? 8'h66 : _GEN_3282; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3284 = 8'hd4 == _t_T_26[15:8] ? 8'h48 : _GEN_3283; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3285 = 8'hd5 == _t_T_26[15:8] ? 8'h3 : _GEN_3284; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3286 = 8'hd6 == _t_T_26[15:8] ? 8'hf6 : _GEN_3285; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3287 = 8'hd7 == _t_T_26[15:8] ? 8'he : _GEN_3286; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3288 = 8'hd8 == _t_T_26[15:8] ? 8'h61 : _GEN_3287; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3289 = 8'hd9 == _t_T_26[15:8] ? 8'h35 : _GEN_3288; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3290 = 8'hda == _t_T_26[15:8] ? 8'h57 : _GEN_3289; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3291 = 8'hdb == _t_T_26[15:8] ? 8'hb9 : _GEN_3290; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3292 = 8'hdc == _t_T_26[15:8] ? 8'h86 : _GEN_3291; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3293 = 8'hdd == _t_T_26[15:8] ? 8'hc1 : _GEN_3292; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3294 = 8'hde == _t_T_26[15:8] ? 8'h1d : _GEN_3293; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3295 = 8'hdf == _t_T_26[15:8] ? 8'h9e : _GEN_3294; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3296 = 8'he0 == _t_T_26[15:8] ? 8'he1 : _GEN_3295; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3297 = 8'he1 == _t_T_26[15:8] ? 8'hf8 : _GEN_3296; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3298 = 8'he2 == _t_T_26[15:8] ? 8'h98 : _GEN_3297; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3299 = 8'he3 == _t_T_26[15:8] ? 8'h11 : _GEN_3298; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3300 = 8'he4 == _t_T_26[15:8] ? 8'h69 : _GEN_3299; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3301 = 8'he5 == _t_T_26[15:8] ? 8'hd9 : _GEN_3300; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3302 = 8'he6 == _t_T_26[15:8] ? 8'h8e : _GEN_3301; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3303 = 8'he7 == _t_T_26[15:8] ? 8'h94 : _GEN_3302; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3304 = 8'he8 == _t_T_26[15:8] ? 8'h9b : _GEN_3303; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3305 = 8'he9 == _t_T_26[15:8] ? 8'h1e : _GEN_3304; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3306 = 8'hea == _t_T_26[15:8] ? 8'h87 : _GEN_3305; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3307 = 8'heb == _t_T_26[15:8] ? 8'he9 : _GEN_3306; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3308 = 8'hec == _t_T_26[15:8] ? 8'hce : _GEN_3307; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3309 = 8'hed == _t_T_26[15:8] ? 8'h55 : _GEN_3308; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3310 = 8'hee == _t_T_26[15:8] ? 8'h28 : _GEN_3309; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3311 = 8'hef == _t_T_26[15:8] ? 8'hdf : _GEN_3310; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3312 = 8'hf0 == _t_T_26[15:8] ? 8'h8c : _GEN_3311; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3313 = 8'hf1 == _t_T_26[15:8] ? 8'ha1 : _GEN_3312; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3314 = 8'hf2 == _t_T_26[15:8] ? 8'h89 : _GEN_3313; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3315 = 8'hf3 == _t_T_26[15:8] ? 8'hd : _GEN_3314; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3316 = 8'hf4 == _t_T_26[15:8] ? 8'hbf : _GEN_3315; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3317 = 8'hf5 == _t_T_26[15:8] ? 8'he6 : _GEN_3316; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3318 = 8'hf6 == _t_T_26[15:8] ? 8'h42 : _GEN_3317; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3319 = 8'hf7 == _t_T_26[15:8] ? 8'h68 : _GEN_3318; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3320 = 8'hf8 == _t_T_26[15:8] ? 8'h41 : _GEN_3319; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3321 = 8'hf9 == _t_T_26[15:8] ? 8'h99 : _GEN_3320; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3322 = 8'hfa == _t_T_26[15:8] ? 8'h2d : _GEN_3321; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3323 = 8'hfb == _t_T_26[15:8] ? 8'hf : _GEN_3322; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3324 = 8'hfc == _t_T_26[15:8] ? 8'hb0 : _GEN_3323; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3325 = 8'hfd == _t_T_26[15:8] ? 8'h54 : _GEN_3324; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3326 = 8'hfe == _t_T_26[15:8] ? 8'hbb : _GEN_3325; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3327 = 8'hff == _t_T_26[15:8] ? 8'h16 : _GEN_3326; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3329 = 8'h1 == _t_T_26[7:0] ? 8'h7c : 8'h63; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3330 = 8'h2 == _t_T_26[7:0] ? 8'h77 : _GEN_3329; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3331 = 8'h3 == _t_T_26[7:0] ? 8'h7b : _GEN_3330; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3332 = 8'h4 == _t_T_26[7:0] ? 8'hf2 : _GEN_3331; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3333 = 8'h5 == _t_T_26[7:0] ? 8'h6b : _GEN_3332; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3334 = 8'h6 == _t_T_26[7:0] ? 8'h6f : _GEN_3333; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3335 = 8'h7 == _t_T_26[7:0] ? 8'hc5 : _GEN_3334; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3336 = 8'h8 == _t_T_26[7:0] ? 8'h30 : _GEN_3335; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3337 = 8'h9 == _t_T_26[7:0] ? 8'h1 : _GEN_3336; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3338 = 8'ha == _t_T_26[7:0] ? 8'h67 : _GEN_3337; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3339 = 8'hb == _t_T_26[7:0] ? 8'h2b : _GEN_3338; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3340 = 8'hc == _t_T_26[7:0] ? 8'hfe : _GEN_3339; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3341 = 8'hd == _t_T_26[7:0] ? 8'hd7 : _GEN_3340; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3342 = 8'he == _t_T_26[7:0] ? 8'hab : _GEN_3341; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3343 = 8'hf == _t_T_26[7:0] ? 8'h76 : _GEN_3342; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3344 = 8'h10 == _t_T_26[7:0] ? 8'hca : _GEN_3343; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3345 = 8'h11 == _t_T_26[7:0] ? 8'h82 : _GEN_3344; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3346 = 8'h12 == _t_T_26[7:0] ? 8'hc9 : _GEN_3345; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3347 = 8'h13 == _t_T_26[7:0] ? 8'h7d : _GEN_3346; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3348 = 8'h14 == _t_T_26[7:0] ? 8'hfa : _GEN_3347; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3349 = 8'h15 == _t_T_26[7:0] ? 8'h59 : _GEN_3348; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3350 = 8'h16 == _t_T_26[7:0] ? 8'h47 : _GEN_3349; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3351 = 8'h17 == _t_T_26[7:0] ? 8'hf0 : _GEN_3350; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3352 = 8'h18 == _t_T_26[7:0] ? 8'had : _GEN_3351; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3353 = 8'h19 == _t_T_26[7:0] ? 8'hd4 : _GEN_3352; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3354 = 8'h1a == _t_T_26[7:0] ? 8'ha2 : _GEN_3353; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3355 = 8'h1b == _t_T_26[7:0] ? 8'haf : _GEN_3354; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3356 = 8'h1c == _t_T_26[7:0] ? 8'h9c : _GEN_3355; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3357 = 8'h1d == _t_T_26[7:0] ? 8'ha4 : _GEN_3356; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3358 = 8'h1e == _t_T_26[7:0] ? 8'h72 : _GEN_3357; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3359 = 8'h1f == _t_T_26[7:0] ? 8'hc0 : _GEN_3358; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3360 = 8'h20 == _t_T_26[7:0] ? 8'hb7 : _GEN_3359; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3361 = 8'h21 == _t_T_26[7:0] ? 8'hfd : _GEN_3360; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3362 = 8'h22 == _t_T_26[7:0] ? 8'h93 : _GEN_3361; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3363 = 8'h23 == _t_T_26[7:0] ? 8'h26 : _GEN_3362; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3364 = 8'h24 == _t_T_26[7:0] ? 8'h36 : _GEN_3363; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3365 = 8'h25 == _t_T_26[7:0] ? 8'h3f : _GEN_3364; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3366 = 8'h26 == _t_T_26[7:0] ? 8'hf7 : _GEN_3365; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3367 = 8'h27 == _t_T_26[7:0] ? 8'hcc : _GEN_3366; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3368 = 8'h28 == _t_T_26[7:0] ? 8'h34 : _GEN_3367; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3369 = 8'h29 == _t_T_26[7:0] ? 8'ha5 : _GEN_3368; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3370 = 8'h2a == _t_T_26[7:0] ? 8'he5 : _GEN_3369; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3371 = 8'h2b == _t_T_26[7:0] ? 8'hf1 : _GEN_3370; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3372 = 8'h2c == _t_T_26[7:0] ? 8'h71 : _GEN_3371; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3373 = 8'h2d == _t_T_26[7:0] ? 8'hd8 : _GEN_3372; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3374 = 8'h2e == _t_T_26[7:0] ? 8'h31 : _GEN_3373; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3375 = 8'h2f == _t_T_26[7:0] ? 8'h15 : _GEN_3374; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3376 = 8'h30 == _t_T_26[7:0] ? 8'h4 : _GEN_3375; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3377 = 8'h31 == _t_T_26[7:0] ? 8'hc7 : _GEN_3376; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3378 = 8'h32 == _t_T_26[7:0] ? 8'h23 : _GEN_3377; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3379 = 8'h33 == _t_T_26[7:0] ? 8'hc3 : _GEN_3378; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3380 = 8'h34 == _t_T_26[7:0] ? 8'h18 : _GEN_3379; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3381 = 8'h35 == _t_T_26[7:0] ? 8'h96 : _GEN_3380; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3382 = 8'h36 == _t_T_26[7:0] ? 8'h5 : _GEN_3381; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3383 = 8'h37 == _t_T_26[7:0] ? 8'h9a : _GEN_3382; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3384 = 8'h38 == _t_T_26[7:0] ? 8'h7 : _GEN_3383; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3385 = 8'h39 == _t_T_26[7:0] ? 8'h12 : _GEN_3384; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3386 = 8'h3a == _t_T_26[7:0] ? 8'h80 : _GEN_3385; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3387 = 8'h3b == _t_T_26[7:0] ? 8'he2 : _GEN_3386; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3388 = 8'h3c == _t_T_26[7:0] ? 8'heb : _GEN_3387; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3389 = 8'h3d == _t_T_26[7:0] ? 8'h27 : _GEN_3388; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3390 = 8'h3e == _t_T_26[7:0] ? 8'hb2 : _GEN_3389; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3391 = 8'h3f == _t_T_26[7:0] ? 8'h75 : _GEN_3390; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3392 = 8'h40 == _t_T_26[7:0] ? 8'h9 : _GEN_3391; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3393 = 8'h41 == _t_T_26[7:0] ? 8'h83 : _GEN_3392; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3394 = 8'h42 == _t_T_26[7:0] ? 8'h2c : _GEN_3393; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3395 = 8'h43 == _t_T_26[7:0] ? 8'h1a : _GEN_3394; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3396 = 8'h44 == _t_T_26[7:0] ? 8'h1b : _GEN_3395; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3397 = 8'h45 == _t_T_26[7:0] ? 8'h6e : _GEN_3396; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3398 = 8'h46 == _t_T_26[7:0] ? 8'h5a : _GEN_3397; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3399 = 8'h47 == _t_T_26[7:0] ? 8'ha0 : _GEN_3398; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3400 = 8'h48 == _t_T_26[7:0] ? 8'h52 : _GEN_3399; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3401 = 8'h49 == _t_T_26[7:0] ? 8'h3b : _GEN_3400; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3402 = 8'h4a == _t_T_26[7:0] ? 8'hd6 : _GEN_3401; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3403 = 8'h4b == _t_T_26[7:0] ? 8'hb3 : _GEN_3402; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3404 = 8'h4c == _t_T_26[7:0] ? 8'h29 : _GEN_3403; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3405 = 8'h4d == _t_T_26[7:0] ? 8'he3 : _GEN_3404; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3406 = 8'h4e == _t_T_26[7:0] ? 8'h2f : _GEN_3405; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3407 = 8'h4f == _t_T_26[7:0] ? 8'h84 : _GEN_3406; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3408 = 8'h50 == _t_T_26[7:0] ? 8'h53 : _GEN_3407; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3409 = 8'h51 == _t_T_26[7:0] ? 8'hd1 : _GEN_3408; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3410 = 8'h52 == _t_T_26[7:0] ? 8'h0 : _GEN_3409; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3411 = 8'h53 == _t_T_26[7:0] ? 8'hed : _GEN_3410; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3412 = 8'h54 == _t_T_26[7:0] ? 8'h20 : _GEN_3411; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3413 = 8'h55 == _t_T_26[7:0] ? 8'hfc : _GEN_3412; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3414 = 8'h56 == _t_T_26[7:0] ? 8'hb1 : _GEN_3413; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3415 = 8'h57 == _t_T_26[7:0] ? 8'h5b : _GEN_3414; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3416 = 8'h58 == _t_T_26[7:0] ? 8'h6a : _GEN_3415; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3417 = 8'h59 == _t_T_26[7:0] ? 8'hcb : _GEN_3416; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3418 = 8'h5a == _t_T_26[7:0] ? 8'hbe : _GEN_3417; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3419 = 8'h5b == _t_T_26[7:0] ? 8'h39 : _GEN_3418; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3420 = 8'h5c == _t_T_26[7:0] ? 8'h4a : _GEN_3419; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3421 = 8'h5d == _t_T_26[7:0] ? 8'h4c : _GEN_3420; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3422 = 8'h5e == _t_T_26[7:0] ? 8'h58 : _GEN_3421; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3423 = 8'h5f == _t_T_26[7:0] ? 8'hcf : _GEN_3422; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3424 = 8'h60 == _t_T_26[7:0] ? 8'hd0 : _GEN_3423; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3425 = 8'h61 == _t_T_26[7:0] ? 8'hef : _GEN_3424; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3426 = 8'h62 == _t_T_26[7:0] ? 8'haa : _GEN_3425; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3427 = 8'h63 == _t_T_26[7:0] ? 8'hfb : _GEN_3426; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3428 = 8'h64 == _t_T_26[7:0] ? 8'h43 : _GEN_3427; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3429 = 8'h65 == _t_T_26[7:0] ? 8'h4d : _GEN_3428; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3430 = 8'h66 == _t_T_26[7:0] ? 8'h33 : _GEN_3429; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3431 = 8'h67 == _t_T_26[7:0] ? 8'h85 : _GEN_3430; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3432 = 8'h68 == _t_T_26[7:0] ? 8'h45 : _GEN_3431; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3433 = 8'h69 == _t_T_26[7:0] ? 8'hf9 : _GEN_3432; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3434 = 8'h6a == _t_T_26[7:0] ? 8'h2 : _GEN_3433; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3435 = 8'h6b == _t_T_26[7:0] ? 8'h7f : _GEN_3434; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3436 = 8'h6c == _t_T_26[7:0] ? 8'h50 : _GEN_3435; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3437 = 8'h6d == _t_T_26[7:0] ? 8'h3c : _GEN_3436; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3438 = 8'h6e == _t_T_26[7:0] ? 8'h9f : _GEN_3437; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3439 = 8'h6f == _t_T_26[7:0] ? 8'ha8 : _GEN_3438; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3440 = 8'h70 == _t_T_26[7:0] ? 8'h51 : _GEN_3439; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3441 = 8'h71 == _t_T_26[7:0] ? 8'ha3 : _GEN_3440; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3442 = 8'h72 == _t_T_26[7:0] ? 8'h40 : _GEN_3441; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3443 = 8'h73 == _t_T_26[7:0] ? 8'h8f : _GEN_3442; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3444 = 8'h74 == _t_T_26[7:0] ? 8'h92 : _GEN_3443; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3445 = 8'h75 == _t_T_26[7:0] ? 8'h9d : _GEN_3444; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3446 = 8'h76 == _t_T_26[7:0] ? 8'h38 : _GEN_3445; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3447 = 8'h77 == _t_T_26[7:0] ? 8'hf5 : _GEN_3446; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3448 = 8'h78 == _t_T_26[7:0] ? 8'hbc : _GEN_3447; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3449 = 8'h79 == _t_T_26[7:0] ? 8'hb6 : _GEN_3448; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3450 = 8'h7a == _t_T_26[7:0] ? 8'hda : _GEN_3449; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3451 = 8'h7b == _t_T_26[7:0] ? 8'h21 : _GEN_3450; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3452 = 8'h7c == _t_T_26[7:0] ? 8'h10 : _GEN_3451; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3453 = 8'h7d == _t_T_26[7:0] ? 8'hff : _GEN_3452; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3454 = 8'h7e == _t_T_26[7:0] ? 8'hf3 : _GEN_3453; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3455 = 8'h7f == _t_T_26[7:0] ? 8'hd2 : _GEN_3454; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3456 = 8'h80 == _t_T_26[7:0] ? 8'hcd : _GEN_3455; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3457 = 8'h81 == _t_T_26[7:0] ? 8'hc : _GEN_3456; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3458 = 8'h82 == _t_T_26[7:0] ? 8'h13 : _GEN_3457; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3459 = 8'h83 == _t_T_26[7:0] ? 8'hec : _GEN_3458; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3460 = 8'h84 == _t_T_26[7:0] ? 8'h5f : _GEN_3459; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3461 = 8'h85 == _t_T_26[7:0] ? 8'h97 : _GEN_3460; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3462 = 8'h86 == _t_T_26[7:0] ? 8'h44 : _GEN_3461; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3463 = 8'h87 == _t_T_26[7:0] ? 8'h17 : _GEN_3462; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3464 = 8'h88 == _t_T_26[7:0] ? 8'hc4 : _GEN_3463; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3465 = 8'h89 == _t_T_26[7:0] ? 8'ha7 : _GEN_3464; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3466 = 8'h8a == _t_T_26[7:0] ? 8'h7e : _GEN_3465; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3467 = 8'h8b == _t_T_26[7:0] ? 8'h3d : _GEN_3466; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3468 = 8'h8c == _t_T_26[7:0] ? 8'h64 : _GEN_3467; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3469 = 8'h8d == _t_T_26[7:0] ? 8'h5d : _GEN_3468; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3470 = 8'h8e == _t_T_26[7:0] ? 8'h19 : _GEN_3469; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3471 = 8'h8f == _t_T_26[7:0] ? 8'h73 : _GEN_3470; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3472 = 8'h90 == _t_T_26[7:0] ? 8'h60 : _GEN_3471; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3473 = 8'h91 == _t_T_26[7:0] ? 8'h81 : _GEN_3472; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3474 = 8'h92 == _t_T_26[7:0] ? 8'h4f : _GEN_3473; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3475 = 8'h93 == _t_T_26[7:0] ? 8'hdc : _GEN_3474; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3476 = 8'h94 == _t_T_26[7:0] ? 8'h22 : _GEN_3475; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3477 = 8'h95 == _t_T_26[7:0] ? 8'h2a : _GEN_3476; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3478 = 8'h96 == _t_T_26[7:0] ? 8'h90 : _GEN_3477; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3479 = 8'h97 == _t_T_26[7:0] ? 8'h88 : _GEN_3478; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3480 = 8'h98 == _t_T_26[7:0] ? 8'h46 : _GEN_3479; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3481 = 8'h99 == _t_T_26[7:0] ? 8'hee : _GEN_3480; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3482 = 8'h9a == _t_T_26[7:0] ? 8'hb8 : _GEN_3481; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3483 = 8'h9b == _t_T_26[7:0] ? 8'h14 : _GEN_3482; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3484 = 8'h9c == _t_T_26[7:0] ? 8'hde : _GEN_3483; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3485 = 8'h9d == _t_T_26[7:0] ? 8'h5e : _GEN_3484; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3486 = 8'h9e == _t_T_26[7:0] ? 8'hb : _GEN_3485; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3487 = 8'h9f == _t_T_26[7:0] ? 8'hdb : _GEN_3486; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3488 = 8'ha0 == _t_T_26[7:0] ? 8'he0 : _GEN_3487; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3489 = 8'ha1 == _t_T_26[7:0] ? 8'h32 : _GEN_3488; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3490 = 8'ha2 == _t_T_26[7:0] ? 8'h3a : _GEN_3489; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3491 = 8'ha3 == _t_T_26[7:0] ? 8'ha : _GEN_3490; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3492 = 8'ha4 == _t_T_26[7:0] ? 8'h49 : _GEN_3491; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3493 = 8'ha5 == _t_T_26[7:0] ? 8'h6 : _GEN_3492; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3494 = 8'ha6 == _t_T_26[7:0] ? 8'h24 : _GEN_3493; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3495 = 8'ha7 == _t_T_26[7:0] ? 8'h5c : _GEN_3494; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3496 = 8'ha8 == _t_T_26[7:0] ? 8'hc2 : _GEN_3495; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3497 = 8'ha9 == _t_T_26[7:0] ? 8'hd3 : _GEN_3496; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3498 = 8'haa == _t_T_26[7:0] ? 8'hac : _GEN_3497; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3499 = 8'hab == _t_T_26[7:0] ? 8'h62 : _GEN_3498; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3500 = 8'hac == _t_T_26[7:0] ? 8'h91 : _GEN_3499; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3501 = 8'had == _t_T_26[7:0] ? 8'h95 : _GEN_3500; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3502 = 8'hae == _t_T_26[7:0] ? 8'he4 : _GEN_3501; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3503 = 8'haf == _t_T_26[7:0] ? 8'h79 : _GEN_3502; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3504 = 8'hb0 == _t_T_26[7:0] ? 8'he7 : _GEN_3503; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3505 = 8'hb1 == _t_T_26[7:0] ? 8'hc8 : _GEN_3504; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3506 = 8'hb2 == _t_T_26[7:0] ? 8'h37 : _GEN_3505; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3507 = 8'hb3 == _t_T_26[7:0] ? 8'h6d : _GEN_3506; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3508 = 8'hb4 == _t_T_26[7:0] ? 8'h8d : _GEN_3507; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3509 = 8'hb5 == _t_T_26[7:0] ? 8'hd5 : _GEN_3508; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3510 = 8'hb6 == _t_T_26[7:0] ? 8'h4e : _GEN_3509; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3511 = 8'hb7 == _t_T_26[7:0] ? 8'ha9 : _GEN_3510; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3512 = 8'hb8 == _t_T_26[7:0] ? 8'h6c : _GEN_3511; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3513 = 8'hb9 == _t_T_26[7:0] ? 8'h56 : _GEN_3512; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3514 = 8'hba == _t_T_26[7:0] ? 8'hf4 : _GEN_3513; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3515 = 8'hbb == _t_T_26[7:0] ? 8'hea : _GEN_3514; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3516 = 8'hbc == _t_T_26[7:0] ? 8'h65 : _GEN_3515; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3517 = 8'hbd == _t_T_26[7:0] ? 8'h7a : _GEN_3516; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3518 = 8'hbe == _t_T_26[7:0] ? 8'hae : _GEN_3517; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3519 = 8'hbf == _t_T_26[7:0] ? 8'h8 : _GEN_3518; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3520 = 8'hc0 == _t_T_26[7:0] ? 8'hba : _GEN_3519; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3521 = 8'hc1 == _t_T_26[7:0] ? 8'h78 : _GEN_3520; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3522 = 8'hc2 == _t_T_26[7:0] ? 8'h25 : _GEN_3521; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3523 = 8'hc3 == _t_T_26[7:0] ? 8'h2e : _GEN_3522; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3524 = 8'hc4 == _t_T_26[7:0] ? 8'h1c : _GEN_3523; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3525 = 8'hc5 == _t_T_26[7:0] ? 8'ha6 : _GEN_3524; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3526 = 8'hc6 == _t_T_26[7:0] ? 8'hb4 : _GEN_3525; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3527 = 8'hc7 == _t_T_26[7:0] ? 8'hc6 : _GEN_3526; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3528 = 8'hc8 == _t_T_26[7:0] ? 8'he8 : _GEN_3527; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3529 = 8'hc9 == _t_T_26[7:0] ? 8'hdd : _GEN_3528; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3530 = 8'hca == _t_T_26[7:0] ? 8'h74 : _GEN_3529; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3531 = 8'hcb == _t_T_26[7:0] ? 8'h1f : _GEN_3530; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3532 = 8'hcc == _t_T_26[7:0] ? 8'h4b : _GEN_3531; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3533 = 8'hcd == _t_T_26[7:0] ? 8'hbd : _GEN_3532; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3534 = 8'hce == _t_T_26[7:0] ? 8'h8b : _GEN_3533; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3535 = 8'hcf == _t_T_26[7:0] ? 8'h8a : _GEN_3534; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3536 = 8'hd0 == _t_T_26[7:0] ? 8'h70 : _GEN_3535; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3537 = 8'hd1 == _t_T_26[7:0] ? 8'h3e : _GEN_3536; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3538 = 8'hd2 == _t_T_26[7:0] ? 8'hb5 : _GEN_3537; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3539 = 8'hd3 == _t_T_26[7:0] ? 8'h66 : _GEN_3538; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3540 = 8'hd4 == _t_T_26[7:0] ? 8'h48 : _GEN_3539; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3541 = 8'hd5 == _t_T_26[7:0] ? 8'h3 : _GEN_3540; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3542 = 8'hd6 == _t_T_26[7:0] ? 8'hf6 : _GEN_3541; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3543 = 8'hd7 == _t_T_26[7:0] ? 8'he : _GEN_3542; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3544 = 8'hd8 == _t_T_26[7:0] ? 8'h61 : _GEN_3543; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3545 = 8'hd9 == _t_T_26[7:0] ? 8'h35 : _GEN_3544; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3546 = 8'hda == _t_T_26[7:0] ? 8'h57 : _GEN_3545; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3547 = 8'hdb == _t_T_26[7:0] ? 8'hb9 : _GEN_3546; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3548 = 8'hdc == _t_T_26[7:0] ? 8'h86 : _GEN_3547; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3549 = 8'hdd == _t_T_26[7:0] ? 8'hc1 : _GEN_3548; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3550 = 8'hde == _t_T_26[7:0] ? 8'h1d : _GEN_3549; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3551 = 8'hdf == _t_T_26[7:0] ? 8'h9e : _GEN_3550; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3552 = 8'he0 == _t_T_26[7:0] ? 8'he1 : _GEN_3551; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3553 = 8'he1 == _t_T_26[7:0] ? 8'hf8 : _GEN_3552; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3554 = 8'he2 == _t_T_26[7:0] ? 8'h98 : _GEN_3553; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3555 = 8'he3 == _t_T_26[7:0] ? 8'h11 : _GEN_3554; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3556 = 8'he4 == _t_T_26[7:0] ? 8'h69 : _GEN_3555; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3557 = 8'he5 == _t_T_26[7:0] ? 8'hd9 : _GEN_3556; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3558 = 8'he6 == _t_T_26[7:0] ? 8'h8e : _GEN_3557; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3559 = 8'he7 == _t_T_26[7:0] ? 8'h94 : _GEN_3558; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3560 = 8'he8 == _t_T_26[7:0] ? 8'h9b : _GEN_3559; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3561 = 8'he9 == _t_T_26[7:0] ? 8'h1e : _GEN_3560; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3562 = 8'hea == _t_T_26[7:0] ? 8'h87 : _GEN_3561; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3563 = 8'heb == _t_T_26[7:0] ? 8'he9 : _GEN_3562; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3564 = 8'hec == _t_T_26[7:0] ? 8'hce : _GEN_3563; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3565 = 8'hed == _t_T_26[7:0] ? 8'h55 : _GEN_3564; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3566 = 8'hee == _t_T_26[7:0] ? 8'h28 : _GEN_3565; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3567 = 8'hef == _t_T_26[7:0] ? 8'hdf : _GEN_3566; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3568 = 8'hf0 == _t_T_26[7:0] ? 8'h8c : _GEN_3567; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3569 = 8'hf1 == _t_T_26[7:0] ? 8'ha1 : _GEN_3568; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3570 = 8'hf2 == _t_T_26[7:0] ? 8'h89 : _GEN_3569; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3571 = 8'hf3 == _t_T_26[7:0] ? 8'hd : _GEN_3570; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3572 = 8'hf4 == _t_T_26[7:0] ? 8'hbf : _GEN_3571; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3573 = 8'hf5 == _t_T_26[7:0] ? 8'he6 : _GEN_3572; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3574 = 8'hf6 == _t_T_26[7:0] ? 8'h42 : _GEN_3573; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3575 = 8'hf7 == _t_T_26[7:0] ? 8'h68 : _GEN_3574; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3576 = 8'hf8 == _t_T_26[7:0] ? 8'h41 : _GEN_3575; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3577 = 8'hf9 == _t_T_26[7:0] ? 8'h99 : _GEN_3576; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3578 = 8'hfa == _t_T_26[7:0] ? 8'h2d : _GEN_3577; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3579 = 8'hfb == _t_T_26[7:0] ? 8'hf : _GEN_3578; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3580 = 8'hfc == _t_T_26[7:0] ? 8'hb0 : _GEN_3579; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3581 = 8'hfd == _t_T_26[7:0] ? 8'h54 : _GEN_3580; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3582 = 8'hfe == _t_T_26[7:0] ? 8'hbb : _GEN_3581; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3583 = 8'hff == _t_T_26[7:0] ? 8'h16 : _GEN_3582; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3585 = 8'h1 == _t_T_26[31:24] ? 8'h7c : 8'h63; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3586 = 8'h2 == _t_T_26[31:24] ? 8'h77 : _GEN_3585; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3587 = 8'h3 == _t_T_26[31:24] ? 8'h7b : _GEN_3586; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3588 = 8'h4 == _t_T_26[31:24] ? 8'hf2 : _GEN_3587; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3589 = 8'h5 == _t_T_26[31:24] ? 8'h6b : _GEN_3588; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3590 = 8'h6 == _t_T_26[31:24] ? 8'h6f : _GEN_3589; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3591 = 8'h7 == _t_T_26[31:24] ? 8'hc5 : _GEN_3590; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3592 = 8'h8 == _t_T_26[31:24] ? 8'h30 : _GEN_3591; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3593 = 8'h9 == _t_T_26[31:24] ? 8'h1 : _GEN_3592; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3594 = 8'ha == _t_T_26[31:24] ? 8'h67 : _GEN_3593; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3595 = 8'hb == _t_T_26[31:24] ? 8'h2b : _GEN_3594; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3596 = 8'hc == _t_T_26[31:24] ? 8'hfe : _GEN_3595; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3597 = 8'hd == _t_T_26[31:24] ? 8'hd7 : _GEN_3596; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3598 = 8'he == _t_T_26[31:24] ? 8'hab : _GEN_3597; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3599 = 8'hf == _t_T_26[31:24] ? 8'h76 : _GEN_3598; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3600 = 8'h10 == _t_T_26[31:24] ? 8'hca : _GEN_3599; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3601 = 8'h11 == _t_T_26[31:24] ? 8'h82 : _GEN_3600; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3602 = 8'h12 == _t_T_26[31:24] ? 8'hc9 : _GEN_3601; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3603 = 8'h13 == _t_T_26[31:24] ? 8'h7d : _GEN_3602; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3604 = 8'h14 == _t_T_26[31:24] ? 8'hfa : _GEN_3603; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3605 = 8'h15 == _t_T_26[31:24] ? 8'h59 : _GEN_3604; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3606 = 8'h16 == _t_T_26[31:24] ? 8'h47 : _GEN_3605; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3607 = 8'h17 == _t_T_26[31:24] ? 8'hf0 : _GEN_3606; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3608 = 8'h18 == _t_T_26[31:24] ? 8'had : _GEN_3607; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3609 = 8'h19 == _t_T_26[31:24] ? 8'hd4 : _GEN_3608; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3610 = 8'h1a == _t_T_26[31:24] ? 8'ha2 : _GEN_3609; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3611 = 8'h1b == _t_T_26[31:24] ? 8'haf : _GEN_3610; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3612 = 8'h1c == _t_T_26[31:24] ? 8'h9c : _GEN_3611; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3613 = 8'h1d == _t_T_26[31:24] ? 8'ha4 : _GEN_3612; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3614 = 8'h1e == _t_T_26[31:24] ? 8'h72 : _GEN_3613; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3615 = 8'h1f == _t_T_26[31:24] ? 8'hc0 : _GEN_3614; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3616 = 8'h20 == _t_T_26[31:24] ? 8'hb7 : _GEN_3615; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3617 = 8'h21 == _t_T_26[31:24] ? 8'hfd : _GEN_3616; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3618 = 8'h22 == _t_T_26[31:24] ? 8'h93 : _GEN_3617; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3619 = 8'h23 == _t_T_26[31:24] ? 8'h26 : _GEN_3618; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3620 = 8'h24 == _t_T_26[31:24] ? 8'h36 : _GEN_3619; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3621 = 8'h25 == _t_T_26[31:24] ? 8'h3f : _GEN_3620; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3622 = 8'h26 == _t_T_26[31:24] ? 8'hf7 : _GEN_3621; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3623 = 8'h27 == _t_T_26[31:24] ? 8'hcc : _GEN_3622; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3624 = 8'h28 == _t_T_26[31:24] ? 8'h34 : _GEN_3623; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3625 = 8'h29 == _t_T_26[31:24] ? 8'ha5 : _GEN_3624; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3626 = 8'h2a == _t_T_26[31:24] ? 8'he5 : _GEN_3625; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3627 = 8'h2b == _t_T_26[31:24] ? 8'hf1 : _GEN_3626; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3628 = 8'h2c == _t_T_26[31:24] ? 8'h71 : _GEN_3627; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3629 = 8'h2d == _t_T_26[31:24] ? 8'hd8 : _GEN_3628; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3630 = 8'h2e == _t_T_26[31:24] ? 8'h31 : _GEN_3629; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3631 = 8'h2f == _t_T_26[31:24] ? 8'h15 : _GEN_3630; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3632 = 8'h30 == _t_T_26[31:24] ? 8'h4 : _GEN_3631; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3633 = 8'h31 == _t_T_26[31:24] ? 8'hc7 : _GEN_3632; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3634 = 8'h32 == _t_T_26[31:24] ? 8'h23 : _GEN_3633; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3635 = 8'h33 == _t_T_26[31:24] ? 8'hc3 : _GEN_3634; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3636 = 8'h34 == _t_T_26[31:24] ? 8'h18 : _GEN_3635; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3637 = 8'h35 == _t_T_26[31:24] ? 8'h96 : _GEN_3636; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3638 = 8'h36 == _t_T_26[31:24] ? 8'h5 : _GEN_3637; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3639 = 8'h37 == _t_T_26[31:24] ? 8'h9a : _GEN_3638; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3640 = 8'h38 == _t_T_26[31:24] ? 8'h7 : _GEN_3639; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3641 = 8'h39 == _t_T_26[31:24] ? 8'h12 : _GEN_3640; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3642 = 8'h3a == _t_T_26[31:24] ? 8'h80 : _GEN_3641; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3643 = 8'h3b == _t_T_26[31:24] ? 8'he2 : _GEN_3642; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3644 = 8'h3c == _t_T_26[31:24] ? 8'heb : _GEN_3643; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3645 = 8'h3d == _t_T_26[31:24] ? 8'h27 : _GEN_3644; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3646 = 8'h3e == _t_T_26[31:24] ? 8'hb2 : _GEN_3645; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3647 = 8'h3f == _t_T_26[31:24] ? 8'h75 : _GEN_3646; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3648 = 8'h40 == _t_T_26[31:24] ? 8'h9 : _GEN_3647; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3649 = 8'h41 == _t_T_26[31:24] ? 8'h83 : _GEN_3648; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3650 = 8'h42 == _t_T_26[31:24] ? 8'h2c : _GEN_3649; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3651 = 8'h43 == _t_T_26[31:24] ? 8'h1a : _GEN_3650; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3652 = 8'h44 == _t_T_26[31:24] ? 8'h1b : _GEN_3651; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3653 = 8'h45 == _t_T_26[31:24] ? 8'h6e : _GEN_3652; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3654 = 8'h46 == _t_T_26[31:24] ? 8'h5a : _GEN_3653; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3655 = 8'h47 == _t_T_26[31:24] ? 8'ha0 : _GEN_3654; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3656 = 8'h48 == _t_T_26[31:24] ? 8'h52 : _GEN_3655; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3657 = 8'h49 == _t_T_26[31:24] ? 8'h3b : _GEN_3656; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3658 = 8'h4a == _t_T_26[31:24] ? 8'hd6 : _GEN_3657; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3659 = 8'h4b == _t_T_26[31:24] ? 8'hb3 : _GEN_3658; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3660 = 8'h4c == _t_T_26[31:24] ? 8'h29 : _GEN_3659; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3661 = 8'h4d == _t_T_26[31:24] ? 8'he3 : _GEN_3660; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3662 = 8'h4e == _t_T_26[31:24] ? 8'h2f : _GEN_3661; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3663 = 8'h4f == _t_T_26[31:24] ? 8'h84 : _GEN_3662; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3664 = 8'h50 == _t_T_26[31:24] ? 8'h53 : _GEN_3663; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3665 = 8'h51 == _t_T_26[31:24] ? 8'hd1 : _GEN_3664; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3666 = 8'h52 == _t_T_26[31:24] ? 8'h0 : _GEN_3665; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3667 = 8'h53 == _t_T_26[31:24] ? 8'hed : _GEN_3666; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3668 = 8'h54 == _t_T_26[31:24] ? 8'h20 : _GEN_3667; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3669 = 8'h55 == _t_T_26[31:24] ? 8'hfc : _GEN_3668; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3670 = 8'h56 == _t_T_26[31:24] ? 8'hb1 : _GEN_3669; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3671 = 8'h57 == _t_T_26[31:24] ? 8'h5b : _GEN_3670; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3672 = 8'h58 == _t_T_26[31:24] ? 8'h6a : _GEN_3671; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3673 = 8'h59 == _t_T_26[31:24] ? 8'hcb : _GEN_3672; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3674 = 8'h5a == _t_T_26[31:24] ? 8'hbe : _GEN_3673; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3675 = 8'h5b == _t_T_26[31:24] ? 8'h39 : _GEN_3674; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3676 = 8'h5c == _t_T_26[31:24] ? 8'h4a : _GEN_3675; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3677 = 8'h5d == _t_T_26[31:24] ? 8'h4c : _GEN_3676; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3678 = 8'h5e == _t_T_26[31:24] ? 8'h58 : _GEN_3677; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3679 = 8'h5f == _t_T_26[31:24] ? 8'hcf : _GEN_3678; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3680 = 8'h60 == _t_T_26[31:24] ? 8'hd0 : _GEN_3679; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3681 = 8'h61 == _t_T_26[31:24] ? 8'hef : _GEN_3680; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3682 = 8'h62 == _t_T_26[31:24] ? 8'haa : _GEN_3681; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3683 = 8'h63 == _t_T_26[31:24] ? 8'hfb : _GEN_3682; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3684 = 8'h64 == _t_T_26[31:24] ? 8'h43 : _GEN_3683; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3685 = 8'h65 == _t_T_26[31:24] ? 8'h4d : _GEN_3684; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3686 = 8'h66 == _t_T_26[31:24] ? 8'h33 : _GEN_3685; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3687 = 8'h67 == _t_T_26[31:24] ? 8'h85 : _GEN_3686; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3688 = 8'h68 == _t_T_26[31:24] ? 8'h45 : _GEN_3687; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3689 = 8'h69 == _t_T_26[31:24] ? 8'hf9 : _GEN_3688; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3690 = 8'h6a == _t_T_26[31:24] ? 8'h2 : _GEN_3689; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3691 = 8'h6b == _t_T_26[31:24] ? 8'h7f : _GEN_3690; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3692 = 8'h6c == _t_T_26[31:24] ? 8'h50 : _GEN_3691; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3693 = 8'h6d == _t_T_26[31:24] ? 8'h3c : _GEN_3692; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3694 = 8'h6e == _t_T_26[31:24] ? 8'h9f : _GEN_3693; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3695 = 8'h6f == _t_T_26[31:24] ? 8'ha8 : _GEN_3694; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3696 = 8'h70 == _t_T_26[31:24] ? 8'h51 : _GEN_3695; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3697 = 8'h71 == _t_T_26[31:24] ? 8'ha3 : _GEN_3696; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3698 = 8'h72 == _t_T_26[31:24] ? 8'h40 : _GEN_3697; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3699 = 8'h73 == _t_T_26[31:24] ? 8'h8f : _GEN_3698; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3700 = 8'h74 == _t_T_26[31:24] ? 8'h92 : _GEN_3699; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3701 = 8'h75 == _t_T_26[31:24] ? 8'h9d : _GEN_3700; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3702 = 8'h76 == _t_T_26[31:24] ? 8'h38 : _GEN_3701; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3703 = 8'h77 == _t_T_26[31:24] ? 8'hf5 : _GEN_3702; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3704 = 8'h78 == _t_T_26[31:24] ? 8'hbc : _GEN_3703; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3705 = 8'h79 == _t_T_26[31:24] ? 8'hb6 : _GEN_3704; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3706 = 8'h7a == _t_T_26[31:24] ? 8'hda : _GEN_3705; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3707 = 8'h7b == _t_T_26[31:24] ? 8'h21 : _GEN_3706; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3708 = 8'h7c == _t_T_26[31:24] ? 8'h10 : _GEN_3707; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3709 = 8'h7d == _t_T_26[31:24] ? 8'hff : _GEN_3708; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3710 = 8'h7e == _t_T_26[31:24] ? 8'hf3 : _GEN_3709; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3711 = 8'h7f == _t_T_26[31:24] ? 8'hd2 : _GEN_3710; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3712 = 8'h80 == _t_T_26[31:24] ? 8'hcd : _GEN_3711; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3713 = 8'h81 == _t_T_26[31:24] ? 8'hc : _GEN_3712; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3714 = 8'h82 == _t_T_26[31:24] ? 8'h13 : _GEN_3713; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3715 = 8'h83 == _t_T_26[31:24] ? 8'hec : _GEN_3714; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3716 = 8'h84 == _t_T_26[31:24] ? 8'h5f : _GEN_3715; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3717 = 8'h85 == _t_T_26[31:24] ? 8'h97 : _GEN_3716; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3718 = 8'h86 == _t_T_26[31:24] ? 8'h44 : _GEN_3717; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3719 = 8'h87 == _t_T_26[31:24] ? 8'h17 : _GEN_3718; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3720 = 8'h88 == _t_T_26[31:24] ? 8'hc4 : _GEN_3719; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3721 = 8'h89 == _t_T_26[31:24] ? 8'ha7 : _GEN_3720; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3722 = 8'h8a == _t_T_26[31:24] ? 8'h7e : _GEN_3721; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3723 = 8'h8b == _t_T_26[31:24] ? 8'h3d : _GEN_3722; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3724 = 8'h8c == _t_T_26[31:24] ? 8'h64 : _GEN_3723; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3725 = 8'h8d == _t_T_26[31:24] ? 8'h5d : _GEN_3724; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3726 = 8'h8e == _t_T_26[31:24] ? 8'h19 : _GEN_3725; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3727 = 8'h8f == _t_T_26[31:24] ? 8'h73 : _GEN_3726; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3728 = 8'h90 == _t_T_26[31:24] ? 8'h60 : _GEN_3727; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3729 = 8'h91 == _t_T_26[31:24] ? 8'h81 : _GEN_3728; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3730 = 8'h92 == _t_T_26[31:24] ? 8'h4f : _GEN_3729; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3731 = 8'h93 == _t_T_26[31:24] ? 8'hdc : _GEN_3730; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3732 = 8'h94 == _t_T_26[31:24] ? 8'h22 : _GEN_3731; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3733 = 8'h95 == _t_T_26[31:24] ? 8'h2a : _GEN_3732; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3734 = 8'h96 == _t_T_26[31:24] ? 8'h90 : _GEN_3733; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3735 = 8'h97 == _t_T_26[31:24] ? 8'h88 : _GEN_3734; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3736 = 8'h98 == _t_T_26[31:24] ? 8'h46 : _GEN_3735; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3737 = 8'h99 == _t_T_26[31:24] ? 8'hee : _GEN_3736; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3738 = 8'h9a == _t_T_26[31:24] ? 8'hb8 : _GEN_3737; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3739 = 8'h9b == _t_T_26[31:24] ? 8'h14 : _GEN_3738; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3740 = 8'h9c == _t_T_26[31:24] ? 8'hde : _GEN_3739; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3741 = 8'h9d == _t_T_26[31:24] ? 8'h5e : _GEN_3740; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3742 = 8'h9e == _t_T_26[31:24] ? 8'hb : _GEN_3741; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3743 = 8'h9f == _t_T_26[31:24] ? 8'hdb : _GEN_3742; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3744 = 8'ha0 == _t_T_26[31:24] ? 8'he0 : _GEN_3743; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3745 = 8'ha1 == _t_T_26[31:24] ? 8'h32 : _GEN_3744; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3746 = 8'ha2 == _t_T_26[31:24] ? 8'h3a : _GEN_3745; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3747 = 8'ha3 == _t_T_26[31:24] ? 8'ha : _GEN_3746; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3748 = 8'ha4 == _t_T_26[31:24] ? 8'h49 : _GEN_3747; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3749 = 8'ha5 == _t_T_26[31:24] ? 8'h6 : _GEN_3748; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3750 = 8'ha6 == _t_T_26[31:24] ? 8'h24 : _GEN_3749; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3751 = 8'ha7 == _t_T_26[31:24] ? 8'h5c : _GEN_3750; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3752 = 8'ha8 == _t_T_26[31:24] ? 8'hc2 : _GEN_3751; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3753 = 8'ha9 == _t_T_26[31:24] ? 8'hd3 : _GEN_3752; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3754 = 8'haa == _t_T_26[31:24] ? 8'hac : _GEN_3753; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3755 = 8'hab == _t_T_26[31:24] ? 8'h62 : _GEN_3754; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3756 = 8'hac == _t_T_26[31:24] ? 8'h91 : _GEN_3755; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3757 = 8'had == _t_T_26[31:24] ? 8'h95 : _GEN_3756; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3758 = 8'hae == _t_T_26[31:24] ? 8'he4 : _GEN_3757; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3759 = 8'haf == _t_T_26[31:24] ? 8'h79 : _GEN_3758; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3760 = 8'hb0 == _t_T_26[31:24] ? 8'he7 : _GEN_3759; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3761 = 8'hb1 == _t_T_26[31:24] ? 8'hc8 : _GEN_3760; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3762 = 8'hb2 == _t_T_26[31:24] ? 8'h37 : _GEN_3761; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3763 = 8'hb3 == _t_T_26[31:24] ? 8'h6d : _GEN_3762; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3764 = 8'hb4 == _t_T_26[31:24] ? 8'h8d : _GEN_3763; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3765 = 8'hb5 == _t_T_26[31:24] ? 8'hd5 : _GEN_3764; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3766 = 8'hb6 == _t_T_26[31:24] ? 8'h4e : _GEN_3765; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3767 = 8'hb7 == _t_T_26[31:24] ? 8'ha9 : _GEN_3766; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3768 = 8'hb8 == _t_T_26[31:24] ? 8'h6c : _GEN_3767; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3769 = 8'hb9 == _t_T_26[31:24] ? 8'h56 : _GEN_3768; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3770 = 8'hba == _t_T_26[31:24] ? 8'hf4 : _GEN_3769; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3771 = 8'hbb == _t_T_26[31:24] ? 8'hea : _GEN_3770; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3772 = 8'hbc == _t_T_26[31:24] ? 8'h65 : _GEN_3771; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3773 = 8'hbd == _t_T_26[31:24] ? 8'h7a : _GEN_3772; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3774 = 8'hbe == _t_T_26[31:24] ? 8'hae : _GEN_3773; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3775 = 8'hbf == _t_T_26[31:24] ? 8'h8 : _GEN_3774; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3776 = 8'hc0 == _t_T_26[31:24] ? 8'hba : _GEN_3775; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3777 = 8'hc1 == _t_T_26[31:24] ? 8'h78 : _GEN_3776; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3778 = 8'hc2 == _t_T_26[31:24] ? 8'h25 : _GEN_3777; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3779 = 8'hc3 == _t_T_26[31:24] ? 8'h2e : _GEN_3778; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3780 = 8'hc4 == _t_T_26[31:24] ? 8'h1c : _GEN_3779; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3781 = 8'hc5 == _t_T_26[31:24] ? 8'ha6 : _GEN_3780; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3782 = 8'hc6 == _t_T_26[31:24] ? 8'hb4 : _GEN_3781; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3783 = 8'hc7 == _t_T_26[31:24] ? 8'hc6 : _GEN_3782; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3784 = 8'hc8 == _t_T_26[31:24] ? 8'he8 : _GEN_3783; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3785 = 8'hc9 == _t_T_26[31:24] ? 8'hdd : _GEN_3784; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3786 = 8'hca == _t_T_26[31:24] ? 8'h74 : _GEN_3785; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3787 = 8'hcb == _t_T_26[31:24] ? 8'h1f : _GEN_3786; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3788 = 8'hcc == _t_T_26[31:24] ? 8'h4b : _GEN_3787; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3789 = 8'hcd == _t_T_26[31:24] ? 8'hbd : _GEN_3788; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3790 = 8'hce == _t_T_26[31:24] ? 8'h8b : _GEN_3789; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3791 = 8'hcf == _t_T_26[31:24] ? 8'h8a : _GEN_3790; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3792 = 8'hd0 == _t_T_26[31:24] ? 8'h70 : _GEN_3791; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3793 = 8'hd1 == _t_T_26[31:24] ? 8'h3e : _GEN_3792; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3794 = 8'hd2 == _t_T_26[31:24] ? 8'hb5 : _GEN_3793; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3795 = 8'hd3 == _t_T_26[31:24] ? 8'h66 : _GEN_3794; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3796 = 8'hd4 == _t_T_26[31:24] ? 8'h48 : _GEN_3795; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3797 = 8'hd5 == _t_T_26[31:24] ? 8'h3 : _GEN_3796; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3798 = 8'hd6 == _t_T_26[31:24] ? 8'hf6 : _GEN_3797; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3799 = 8'hd7 == _t_T_26[31:24] ? 8'he : _GEN_3798; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3800 = 8'hd8 == _t_T_26[31:24] ? 8'h61 : _GEN_3799; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3801 = 8'hd9 == _t_T_26[31:24] ? 8'h35 : _GEN_3800; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3802 = 8'hda == _t_T_26[31:24] ? 8'h57 : _GEN_3801; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3803 = 8'hdb == _t_T_26[31:24] ? 8'hb9 : _GEN_3802; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3804 = 8'hdc == _t_T_26[31:24] ? 8'h86 : _GEN_3803; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3805 = 8'hdd == _t_T_26[31:24] ? 8'hc1 : _GEN_3804; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3806 = 8'hde == _t_T_26[31:24] ? 8'h1d : _GEN_3805; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3807 = 8'hdf == _t_T_26[31:24] ? 8'h9e : _GEN_3806; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3808 = 8'he0 == _t_T_26[31:24] ? 8'he1 : _GEN_3807; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3809 = 8'he1 == _t_T_26[31:24] ? 8'hf8 : _GEN_3808; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3810 = 8'he2 == _t_T_26[31:24] ? 8'h98 : _GEN_3809; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3811 = 8'he3 == _t_T_26[31:24] ? 8'h11 : _GEN_3810; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3812 = 8'he4 == _t_T_26[31:24] ? 8'h69 : _GEN_3811; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3813 = 8'he5 == _t_T_26[31:24] ? 8'hd9 : _GEN_3812; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3814 = 8'he6 == _t_T_26[31:24] ? 8'h8e : _GEN_3813; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3815 = 8'he7 == _t_T_26[31:24] ? 8'h94 : _GEN_3814; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3816 = 8'he8 == _t_T_26[31:24] ? 8'h9b : _GEN_3815; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3817 = 8'he9 == _t_T_26[31:24] ? 8'h1e : _GEN_3816; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3818 = 8'hea == _t_T_26[31:24] ? 8'h87 : _GEN_3817; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3819 = 8'heb == _t_T_26[31:24] ? 8'he9 : _GEN_3818; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3820 = 8'hec == _t_T_26[31:24] ? 8'hce : _GEN_3819; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3821 = 8'hed == _t_T_26[31:24] ? 8'h55 : _GEN_3820; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3822 = 8'hee == _t_T_26[31:24] ? 8'h28 : _GEN_3821; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3823 = 8'hef == _t_T_26[31:24] ? 8'hdf : _GEN_3822; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3824 = 8'hf0 == _t_T_26[31:24] ? 8'h8c : _GEN_3823; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3825 = 8'hf1 == _t_T_26[31:24] ? 8'ha1 : _GEN_3824; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3826 = 8'hf2 == _t_T_26[31:24] ? 8'h89 : _GEN_3825; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3827 = 8'hf3 == _t_T_26[31:24] ? 8'hd : _GEN_3826; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3828 = 8'hf4 == _t_T_26[31:24] ? 8'hbf : _GEN_3827; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3829 = 8'hf5 == _t_T_26[31:24] ? 8'he6 : _GEN_3828; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3830 = 8'hf6 == _t_T_26[31:24] ? 8'h42 : _GEN_3829; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3831 = 8'hf7 == _t_T_26[31:24] ? 8'h68 : _GEN_3830; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3832 = 8'hf8 == _t_T_26[31:24] ? 8'h41 : _GEN_3831; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3833 = 8'hf9 == _t_T_26[31:24] ? 8'h99 : _GEN_3832; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3834 = 8'hfa == _t_T_26[31:24] ? 8'h2d : _GEN_3833; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3835 = 8'hfb == _t_T_26[31:24] ? 8'hf : _GEN_3834; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3836 = 8'hfc == _t_T_26[31:24] ? 8'hb0 : _GEN_3835; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3837 = 8'hfd == _t_T_26[31:24] ? 8'h54 : _GEN_3836; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3838 = 8'hfe == _t_T_26[31:24] ? 8'hbb : _GEN_3837; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3839 = 8'hff == _t_T_26[31:24] ? 8'h16 : _GEN_3838; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3841 = 8'h1 == _t_T_26[23:16] ? 8'h7c : 8'h63; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3842 = 8'h2 == _t_T_26[23:16] ? 8'h77 : _GEN_3841; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3843 = 8'h3 == _t_T_26[23:16] ? 8'h7b : _GEN_3842; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3844 = 8'h4 == _t_T_26[23:16] ? 8'hf2 : _GEN_3843; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3845 = 8'h5 == _t_T_26[23:16] ? 8'h6b : _GEN_3844; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3846 = 8'h6 == _t_T_26[23:16] ? 8'h6f : _GEN_3845; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3847 = 8'h7 == _t_T_26[23:16] ? 8'hc5 : _GEN_3846; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3848 = 8'h8 == _t_T_26[23:16] ? 8'h30 : _GEN_3847; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3849 = 8'h9 == _t_T_26[23:16] ? 8'h1 : _GEN_3848; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3850 = 8'ha == _t_T_26[23:16] ? 8'h67 : _GEN_3849; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3851 = 8'hb == _t_T_26[23:16] ? 8'h2b : _GEN_3850; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3852 = 8'hc == _t_T_26[23:16] ? 8'hfe : _GEN_3851; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3853 = 8'hd == _t_T_26[23:16] ? 8'hd7 : _GEN_3852; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3854 = 8'he == _t_T_26[23:16] ? 8'hab : _GEN_3853; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3855 = 8'hf == _t_T_26[23:16] ? 8'h76 : _GEN_3854; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3856 = 8'h10 == _t_T_26[23:16] ? 8'hca : _GEN_3855; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3857 = 8'h11 == _t_T_26[23:16] ? 8'h82 : _GEN_3856; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3858 = 8'h12 == _t_T_26[23:16] ? 8'hc9 : _GEN_3857; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3859 = 8'h13 == _t_T_26[23:16] ? 8'h7d : _GEN_3858; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3860 = 8'h14 == _t_T_26[23:16] ? 8'hfa : _GEN_3859; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3861 = 8'h15 == _t_T_26[23:16] ? 8'h59 : _GEN_3860; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3862 = 8'h16 == _t_T_26[23:16] ? 8'h47 : _GEN_3861; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3863 = 8'h17 == _t_T_26[23:16] ? 8'hf0 : _GEN_3862; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3864 = 8'h18 == _t_T_26[23:16] ? 8'had : _GEN_3863; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3865 = 8'h19 == _t_T_26[23:16] ? 8'hd4 : _GEN_3864; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3866 = 8'h1a == _t_T_26[23:16] ? 8'ha2 : _GEN_3865; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3867 = 8'h1b == _t_T_26[23:16] ? 8'haf : _GEN_3866; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3868 = 8'h1c == _t_T_26[23:16] ? 8'h9c : _GEN_3867; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3869 = 8'h1d == _t_T_26[23:16] ? 8'ha4 : _GEN_3868; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3870 = 8'h1e == _t_T_26[23:16] ? 8'h72 : _GEN_3869; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3871 = 8'h1f == _t_T_26[23:16] ? 8'hc0 : _GEN_3870; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3872 = 8'h20 == _t_T_26[23:16] ? 8'hb7 : _GEN_3871; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3873 = 8'h21 == _t_T_26[23:16] ? 8'hfd : _GEN_3872; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3874 = 8'h22 == _t_T_26[23:16] ? 8'h93 : _GEN_3873; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3875 = 8'h23 == _t_T_26[23:16] ? 8'h26 : _GEN_3874; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3876 = 8'h24 == _t_T_26[23:16] ? 8'h36 : _GEN_3875; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3877 = 8'h25 == _t_T_26[23:16] ? 8'h3f : _GEN_3876; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3878 = 8'h26 == _t_T_26[23:16] ? 8'hf7 : _GEN_3877; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3879 = 8'h27 == _t_T_26[23:16] ? 8'hcc : _GEN_3878; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3880 = 8'h28 == _t_T_26[23:16] ? 8'h34 : _GEN_3879; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3881 = 8'h29 == _t_T_26[23:16] ? 8'ha5 : _GEN_3880; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3882 = 8'h2a == _t_T_26[23:16] ? 8'he5 : _GEN_3881; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3883 = 8'h2b == _t_T_26[23:16] ? 8'hf1 : _GEN_3882; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3884 = 8'h2c == _t_T_26[23:16] ? 8'h71 : _GEN_3883; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3885 = 8'h2d == _t_T_26[23:16] ? 8'hd8 : _GEN_3884; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3886 = 8'h2e == _t_T_26[23:16] ? 8'h31 : _GEN_3885; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3887 = 8'h2f == _t_T_26[23:16] ? 8'h15 : _GEN_3886; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3888 = 8'h30 == _t_T_26[23:16] ? 8'h4 : _GEN_3887; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3889 = 8'h31 == _t_T_26[23:16] ? 8'hc7 : _GEN_3888; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3890 = 8'h32 == _t_T_26[23:16] ? 8'h23 : _GEN_3889; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3891 = 8'h33 == _t_T_26[23:16] ? 8'hc3 : _GEN_3890; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3892 = 8'h34 == _t_T_26[23:16] ? 8'h18 : _GEN_3891; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3893 = 8'h35 == _t_T_26[23:16] ? 8'h96 : _GEN_3892; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3894 = 8'h36 == _t_T_26[23:16] ? 8'h5 : _GEN_3893; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3895 = 8'h37 == _t_T_26[23:16] ? 8'h9a : _GEN_3894; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3896 = 8'h38 == _t_T_26[23:16] ? 8'h7 : _GEN_3895; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3897 = 8'h39 == _t_T_26[23:16] ? 8'h12 : _GEN_3896; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3898 = 8'h3a == _t_T_26[23:16] ? 8'h80 : _GEN_3897; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3899 = 8'h3b == _t_T_26[23:16] ? 8'he2 : _GEN_3898; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3900 = 8'h3c == _t_T_26[23:16] ? 8'heb : _GEN_3899; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3901 = 8'h3d == _t_T_26[23:16] ? 8'h27 : _GEN_3900; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3902 = 8'h3e == _t_T_26[23:16] ? 8'hb2 : _GEN_3901; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3903 = 8'h3f == _t_T_26[23:16] ? 8'h75 : _GEN_3902; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3904 = 8'h40 == _t_T_26[23:16] ? 8'h9 : _GEN_3903; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3905 = 8'h41 == _t_T_26[23:16] ? 8'h83 : _GEN_3904; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3906 = 8'h42 == _t_T_26[23:16] ? 8'h2c : _GEN_3905; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3907 = 8'h43 == _t_T_26[23:16] ? 8'h1a : _GEN_3906; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3908 = 8'h44 == _t_T_26[23:16] ? 8'h1b : _GEN_3907; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3909 = 8'h45 == _t_T_26[23:16] ? 8'h6e : _GEN_3908; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3910 = 8'h46 == _t_T_26[23:16] ? 8'h5a : _GEN_3909; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3911 = 8'h47 == _t_T_26[23:16] ? 8'ha0 : _GEN_3910; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3912 = 8'h48 == _t_T_26[23:16] ? 8'h52 : _GEN_3911; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3913 = 8'h49 == _t_T_26[23:16] ? 8'h3b : _GEN_3912; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3914 = 8'h4a == _t_T_26[23:16] ? 8'hd6 : _GEN_3913; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3915 = 8'h4b == _t_T_26[23:16] ? 8'hb3 : _GEN_3914; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3916 = 8'h4c == _t_T_26[23:16] ? 8'h29 : _GEN_3915; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3917 = 8'h4d == _t_T_26[23:16] ? 8'he3 : _GEN_3916; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3918 = 8'h4e == _t_T_26[23:16] ? 8'h2f : _GEN_3917; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3919 = 8'h4f == _t_T_26[23:16] ? 8'h84 : _GEN_3918; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3920 = 8'h50 == _t_T_26[23:16] ? 8'h53 : _GEN_3919; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3921 = 8'h51 == _t_T_26[23:16] ? 8'hd1 : _GEN_3920; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3922 = 8'h52 == _t_T_26[23:16] ? 8'h0 : _GEN_3921; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3923 = 8'h53 == _t_T_26[23:16] ? 8'hed : _GEN_3922; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3924 = 8'h54 == _t_T_26[23:16] ? 8'h20 : _GEN_3923; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3925 = 8'h55 == _t_T_26[23:16] ? 8'hfc : _GEN_3924; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3926 = 8'h56 == _t_T_26[23:16] ? 8'hb1 : _GEN_3925; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3927 = 8'h57 == _t_T_26[23:16] ? 8'h5b : _GEN_3926; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3928 = 8'h58 == _t_T_26[23:16] ? 8'h6a : _GEN_3927; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3929 = 8'h59 == _t_T_26[23:16] ? 8'hcb : _GEN_3928; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3930 = 8'h5a == _t_T_26[23:16] ? 8'hbe : _GEN_3929; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3931 = 8'h5b == _t_T_26[23:16] ? 8'h39 : _GEN_3930; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3932 = 8'h5c == _t_T_26[23:16] ? 8'h4a : _GEN_3931; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3933 = 8'h5d == _t_T_26[23:16] ? 8'h4c : _GEN_3932; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3934 = 8'h5e == _t_T_26[23:16] ? 8'h58 : _GEN_3933; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3935 = 8'h5f == _t_T_26[23:16] ? 8'hcf : _GEN_3934; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3936 = 8'h60 == _t_T_26[23:16] ? 8'hd0 : _GEN_3935; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3937 = 8'h61 == _t_T_26[23:16] ? 8'hef : _GEN_3936; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3938 = 8'h62 == _t_T_26[23:16] ? 8'haa : _GEN_3937; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3939 = 8'h63 == _t_T_26[23:16] ? 8'hfb : _GEN_3938; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3940 = 8'h64 == _t_T_26[23:16] ? 8'h43 : _GEN_3939; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3941 = 8'h65 == _t_T_26[23:16] ? 8'h4d : _GEN_3940; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3942 = 8'h66 == _t_T_26[23:16] ? 8'h33 : _GEN_3941; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3943 = 8'h67 == _t_T_26[23:16] ? 8'h85 : _GEN_3942; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3944 = 8'h68 == _t_T_26[23:16] ? 8'h45 : _GEN_3943; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3945 = 8'h69 == _t_T_26[23:16] ? 8'hf9 : _GEN_3944; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3946 = 8'h6a == _t_T_26[23:16] ? 8'h2 : _GEN_3945; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3947 = 8'h6b == _t_T_26[23:16] ? 8'h7f : _GEN_3946; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3948 = 8'h6c == _t_T_26[23:16] ? 8'h50 : _GEN_3947; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3949 = 8'h6d == _t_T_26[23:16] ? 8'h3c : _GEN_3948; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3950 = 8'h6e == _t_T_26[23:16] ? 8'h9f : _GEN_3949; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3951 = 8'h6f == _t_T_26[23:16] ? 8'ha8 : _GEN_3950; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3952 = 8'h70 == _t_T_26[23:16] ? 8'h51 : _GEN_3951; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3953 = 8'h71 == _t_T_26[23:16] ? 8'ha3 : _GEN_3952; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3954 = 8'h72 == _t_T_26[23:16] ? 8'h40 : _GEN_3953; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3955 = 8'h73 == _t_T_26[23:16] ? 8'h8f : _GEN_3954; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3956 = 8'h74 == _t_T_26[23:16] ? 8'h92 : _GEN_3955; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3957 = 8'h75 == _t_T_26[23:16] ? 8'h9d : _GEN_3956; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3958 = 8'h76 == _t_T_26[23:16] ? 8'h38 : _GEN_3957; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3959 = 8'h77 == _t_T_26[23:16] ? 8'hf5 : _GEN_3958; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3960 = 8'h78 == _t_T_26[23:16] ? 8'hbc : _GEN_3959; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3961 = 8'h79 == _t_T_26[23:16] ? 8'hb6 : _GEN_3960; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3962 = 8'h7a == _t_T_26[23:16] ? 8'hda : _GEN_3961; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3963 = 8'h7b == _t_T_26[23:16] ? 8'h21 : _GEN_3962; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3964 = 8'h7c == _t_T_26[23:16] ? 8'h10 : _GEN_3963; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3965 = 8'h7d == _t_T_26[23:16] ? 8'hff : _GEN_3964; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3966 = 8'h7e == _t_T_26[23:16] ? 8'hf3 : _GEN_3965; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3967 = 8'h7f == _t_T_26[23:16] ? 8'hd2 : _GEN_3966; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3968 = 8'h80 == _t_T_26[23:16] ? 8'hcd : _GEN_3967; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3969 = 8'h81 == _t_T_26[23:16] ? 8'hc : _GEN_3968; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3970 = 8'h82 == _t_T_26[23:16] ? 8'h13 : _GEN_3969; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3971 = 8'h83 == _t_T_26[23:16] ? 8'hec : _GEN_3970; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3972 = 8'h84 == _t_T_26[23:16] ? 8'h5f : _GEN_3971; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3973 = 8'h85 == _t_T_26[23:16] ? 8'h97 : _GEN_3972; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3974 = 8'h86 == _t_T_26[23:16] ? 8'h44 : _GEN_3973; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3975 = 8'h87 == _t_T_26[23:16] ? 8'h17 : _GEN_3974; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3976 = 8'h88 == _t_T_26[23:16] ? 8'hc4 : _GEN_3975; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3977 = 8'h89 == _t_T_26[23:16] ? 8'ha7 : _GEN_3976; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3978 = 8'h8a == _t_T_26[23:16] ? 8'h7e : _GEN_3977; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3979 = 8'h8b == _t_T_26[23:16] ? 8'h3d : _GEN_3978; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3980 = 8'h8c == _t_T_26[23:16] ? 8'h64 : _GEN_3979; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3981 = 8'h8d == _t_T_26[23:16] ? 8'h5d : _GEN_3980; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3982 = 8'h8e == _t_T_26[23:16] ? 8'h19 : _GEN_3981; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3983 = 8'h8f == _t_T_26[23:16] ? 8'h73 : _GEN_3982; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3984 = 8'h90 == _t_T_26[23:16] ? 8'h60 : _GEN_3983; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3985 = 8'h91 == _t_T_26[23:16] ? 8'h81 : _GEN_3984; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3986 = 8'h92 == _t_T_26[23:16] ? 8'h4f : _GEN_3985; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3987 = 8'h93 == _t_T_26[23:16] ? 8'hdc : _GEN_3986; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3988 = 8'h94 == _t_T_26[23:16] ? 8'h22 : _GEN_3987; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3989 = 8'h95 == _t_T_26[23:16] ? 8'h2a : _GEN_3988; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3990 = 8'h96 == _t_T_26[23:16] ? 8'h90 : _GEN_3989; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3991 = 8'h97 == _t_T_26[23:16] ? 8'h88 : _GEN_3990; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3992 = 8'h98 == _t_T_26[23:16] ? 8'h46 : _GEN_3991; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3993 = 8'h99 == _t_T_26[23:16] ? 8'hee : _GEN_3992; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3994 = 8'h9a == _t_T_26[23:16] ? 8'hb8 : _GEN_3993; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3995 = 8'h9b == _t_T_26[23:16] ? 8'h14 : _GEN_3994; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3996 = 8'h9c == _t_T_26[23:16] ? 8'hde : _GEN_3995; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3997 = 8'h9d == _t_T_26[23:16] ? 8'h5e : _GEN_3996; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3998 = 8'h9e == _t_T_26[23:16] ? 8'hb : _GEN_3997; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_3999 = 8'h9f == _t_T_26[23:16] ? 8'hdb : _GEN_3998; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4000 = 8'ha0 == _t_T_26[23:16] ? 8'he0 : _GEN_3999; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4001 = 8'ha1 == _t_T_26[23:16] ? 8'h32 : _GEN_4000; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4002 = 8'ha2 == _t_T_26[23:16] ? 8'h3a : _GEN_4001; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4003 = 8'ha3 == _t_T_26[23:16] ? 8'ha : _GEN_4002; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4004 = 8'ha4 == _t_T_26[23:16] ? 8'h49 : _GEN_4003; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4005 = 8'ha5 == _t_T_26[23:16] ? 8'h6 : _GEN_4004; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4006 = 8'ha6 == _t_T_26[23:16] ? 8'h24 : _GEN_4005; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4007 = 8'ha7 == _t_T_26[23:16] ? 8'h5c : _GEN_4006; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4008 = 8'ha8 == _t_T_26[23:16] ? 8'hc2 : _GEN_4007; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4009 = 8'ha9 == _t_T_26[23:16] ? 8'hd3 : _GEN_4008; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4010 = 8'haa == _t_T_26[23:16] ? 8'hac : _GEN_4009; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4011 = 8'hab == _t_T_26[23:16] ? 8'h62 : _GEN_4010; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4012 = 8'hac == _t_T_26[23:16] ? 8'h91 : _GEN_4011; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4013 = 8'had == _t_T_26[23:16] ? 8'h95 : _GEN_4012; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4014 = 8'hae == _t_T_26[23:16] ? 8'he4 : _GEN_4013; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4015 = 8'haf == _t_T_26[23:16] ? 8'h79 : _GEN_4014; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4016 = 8'hb0 == _t_T_26[23:16] ? 8'he7 : _GEN_4015; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4017 = 8'hb1 == _t_T_26[23:16] ? 8'hc8 : _GEN_4016; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4018 = 8'hb2 == _t_T_26[23:16] ? 8'h37 : _GEN_4017; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4019 = 8'hb3 == _t_T_26[23:16] ? 8'h6d : _GEN_4018; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4020 = 8'hb4 == _t_T_26[23:16] ? 8'h8d : _GEN_4019; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4021 = 8'hb5 == _t_T_26[23:16] ? 8'hd5 : _GEN_4020; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4022 = 8'hb6 == _t_T_26[23:16] ? 8'h4e : _GEN_4021; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4023 = 8'hb7 == _t_T_26[23:16] ? 8'ha9 : _GEN_4022; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4024 = 8'hb8 == _t_T_26[23:16] ? 8'h6c : _GEN_4023; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4025 = 8'hb9 == _t_T_26[23:16] ? 8'h56 : _GEN_4024; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4026 = 8'hba == _t_T_26[23:16] ? 8'hf4 : _GEN_4025; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4027 = 8'hbb == _t_T_26[23:16] ? 8'hea : _GEN_4026; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4028 = 8'hbc == _t_T_26[23:16] ? 8'h65 : _GEN_4027; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4029 = 8'hbd == _t_T_26[23:16] ? 8'h7a : _GEN_4028; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4030 = 8'hbe == _t_T_26[23:16] ? 8'hae : _GEN_4029; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4031 = 8'hbf == _t_T_26[23:16] ? 8'h8 : _GEN_4030; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4032 = 8'hc0 == _t_T_26[23:16] ? 8'hba : _GEN_4031; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4033 = 8'hc1 == _t_T_26[23:16] ? 8'h78 : _GEN_4032; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4034 = 8'hc2 == _t_T_26[23:16] ? 8'h25 : _GEN_4033; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4035 = 8'hc3 == _t_T_26[23:16] ? 8'h2e : _GEN_4034; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4036 = 8'hc4 == _t_T_26[23:16] ? 8'h1c : _GEN_4035; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4037 = 8'hc5 == _t_T_26[23:16] ? 8'ha6 : _GEN_4036; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4038 = 8'hc6 == _t_T_26[23:16] ? 8'hb4 : _GEN_4037; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4039 = 8'hc7 == _t_T_26[23:16] ? 8'hc6 : _GEN_4038; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4040 = 8'hc8 == _t_T_26[23:16] ? 8'he8 : _GEN_4039; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4041 = 8'hc9 == _t_T_26[23:16] ? 8'hdd : _GEN_4040; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4042 = 8'hca == _t_T_26[23:16] ? 8'h74 : _GEN_4041; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4043 = 8'hcb == _t_T_26[23:16] ? 8'h1f : _GEN_4042; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4044 = 8'hcc == _t_T_26[23:16] ? 8'h4b : _GEN_4043; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4045 = 8'hcd == _t_T_26[23:16] ? 8'hbd : _GEN_4044; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4046 = 8'hce == _t_T_26[23:16] ? 8'h8b : _GEN_4045; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4047 = 8'hcf == _t_T_26[23:16] ? 8'h8a : _GEN_4046; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4048 = 8'hd0 == _t_T_26[23:16] ? 8'h70 : _GEN_4047; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4049 = 8'hd1 == _t_T_26[23:16] ? 8'h3e : _GEN_4048; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4050 = 8'hd2 == _t_T_26[23:16] ? 8'hb5 : _GEN_4049; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4051 = 8'hd3 == _t_T_26[23:16] ? 8'h66 : _GEN_4050; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4052 = 8'hd4 == _t_T_26[23:16] ? 8'h48 : _GEN_4051; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4053 = 8'hd5 == _t_T_26[23:16] ? 8'h3 : _GEN_4052; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4054 = 8'hd6 == _t_T_26[23:16] ? 8'hf6 : _GEN_4053; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4055 = 8'hd7 == _t_T_26[23:16] ? 8'he : _GEN_4054; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4056 = 8'hd8 == _t_T_26[23:16] ? 8'h61 : _GEN_4055; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4057 = 8'hd9 == _t_T_26[23:16] ? 8'h35 : _GEN_4056; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4058 = 8'hda == _t_T_26[23:16] ? 8'h57 : _GEN_4057; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4059 = 8'hdb == _t_T_26[23:16] ? 8'hb9 : _GEN_4058; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4060 = 8'hdc == _t_T_26[23:16] ? 8'h86 : _GEN_4059; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4061 = 8'hdd == _t_T_26[23:16] ? 8'hc1 : _GEN_4060; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4062 = 8'hde == _t_T_26[23:16] ? 8'h1d : _GEN_4061; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4063 = 8'hdf == _t_T_26[23:16] ? 8'h9e : _GEN_4062; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4064 = 8'he0 == _t_T_26[23:16] ? 8'he1 : _GEN_4063; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4065 = 8'he1 == _t_T_26[23:16] ? 8'hf8 : _GEN_4064; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4066 = 8'he2 == _t_T_26[23:16] ? 8'h98 : _GEN_4065; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4067 = 8'he3 == _t_T_26[23:16] ? 8'h11 : _GEN_4066; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4068 = 8'he4 == _t_T_26[23:16] ? 8'h69 : _GEN_4067; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4069 = 8'he5 == _t_T_26[23:16] ? 8'hd9 : _GEN_4068; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4070 = 8'he6 == _t_T_26[23:16] ? 8'h8e : _GEN_4069; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4071 = 8'he7 == _t_T_26[23:16] ? 8'h94 : _GEN_4070; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4072 = 8'he8 == _t_T_26[23:16] ? 8'h9b : _GEN_4071; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4073 = 8'he9 == _t_T_26[23:16] ? 8'h1e : _GEN_4072; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4074 = 8'hea == _t_T_26[23:16] ? 8'h87 : _GEN_4073; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4075 = 8'heb == _t_T_26[23:16] ? 8'he9 : _GEN_4074; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4076 = 8'hec == _t_T_26[23:16] ? 8'hce : _GEN_4075; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4077 = 8'hed == _t_T_26[23:16] ? 8'h55 : _GEN_4076; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4078 = 8'hee == _t_T_26[23:16] ? 8'h28 : _GEN_4077; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4079 = 8'hef == _t_T_26[23:16] ? 8'hdf : _GEN_4078; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4080 = 8'hf0 == _t_T_26[23:16] ? 8'h8c : _GEN_4079; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4081 = 8'hf1 == _t_T_26[23:16] ? 8'ha1 : _GEN_4080; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4082 = 8'hf2 == _t_T_26[23:16] ? 8'h89 : _GEN_4081; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4083 = 8'hf3 == _t_T_26[23:16] ? 8'hd : _GEN_4082; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4084 = 8'hf4 == _t_T_26[23:16] ? 8'hbf : _GEN_4083; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4085 = 8'hf5 == _t_T_26[23:16] ? 8'he6 : _GEN_4084; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4086 = 8'hf6 == _t_T_26[23:16] ? 8'h42 : _GEN_4085; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4087 = 8'hf7 == _t_T_26[23:16] ? 8'h68 : _GEN_4086; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4088 = 8'hf8 == _t_T_26[23:16] ? 8'h41 : _GEN_4087; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4089 = 8'hf9 == _t_T_26[23:16] ? 8'h99 : _GEN_4088; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4090 = 8'hfa == _t_T_26[23:16] ? 8'h2d : _GEN_4089; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4091 = 8'hfb == _t_T_26[23:16] ? 8'hf : _GEN_4090; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4092 = 8'hfc == _t_T_26[23:16] ? 8'hb0 : _GEN_4091; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4093 = 8'hfd == _t_T_26[23:16] ? 8'h54 : _GEN_4092; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4094 = 8'hfe == _t_T_26[23:16] ? 8'hbb : _GEN_4093; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4095 = 8'hff == _t_T_26[23:16] ? 8'h16 : _GEN_4094; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [31:0] _t_T_31 = {_GEN_3839,_GEN_4095,_GEN_3327,_GEN_3583}; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:8]
  wire [31:0] t_3 = _t_T_31 ^ 32'h8000000; // @[src/main/scala/crypto/aes/KeySchedule.scala 59:32]
  wire [31:0] w_16 = w_12 ^ t_3; // @[src/main/scala/crypto/aes/KeySchedule.scala 63:21]
  wire [31:0] w_17 = w_13 ^ w_16; // @[src/main/scala/crypto/aes/KeySchedule.scala 63:21]
  wire [31:0] w_18 = w_14 ^ w_17; // @[src/main/scala/crypto/aes/KeySchedule.scala 63:21]
  wire [31:0] w_19 = w_15 ^ w_18; // @[src/main/scala/crypto/aes/KeySchedule.scala 63:21]
  wire [31:0] _t_T_34 = {w_19[23:0],w_19[31:24]}; // @[src/main/scala/crypto/aes/KeySchedule.scala 23:43]
  wire [7:0] _GEN_4097 = 8'h1 == _t_T_34[15:8] ? 8'h7c : 8'h63; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4098 = 8'h2 == _t_T_34[15:8] ? 8'h77 : _GEN_4097; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4099 = 8'h3 == _t_T_34[15:8] ? 8'h7b : _GEN_4098; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4100 = 8'h4 == _t_T_34[15:8] ? 8'hf2 : _GEN_4099; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4101 = 8'h5 == _t_T_34[15:8] ? 8'h6b : _GEN_4100; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4102 = 8'h6 == _t_T_34[15:8] ? 8'h6f : _GEN_4101; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4103 = 8'h7 == _t_T_34[15:8] ? 8'hc5 : _GEN_4102; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4104 = 8'h8 == _t_T_34[15:8] ? 8'h30 : _GEN_4103; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4105 = 8'h9 == _t_T_34[15:8] ? 8'h1 : _GEN_4104; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4106 = 8'ha == _t_T_34[15:8] ? 8'h67 : _GEN_4105; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4107 = 8'hb == _t_T_34[15:8] ? 8'h2b : _GEN_4106; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4108 = 8'hc == _t_T_34[15:8] ? 8'hfe : _GEN_4107; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4109 = 8'hd == _t_T_34[15:8] ? 8'hd7 : _GEN_4108; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4110 = 8'he == _t_T_34[15:8] ? 8'hab : _GEN_4109; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4111 = 8'hf == _t_T_34[15:8] ? 8'h76 : _GEN_4110; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4112 = 8'h10 == _t_T_34[15:8] ? 8'hca : _GEN_4111; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4113 = 8'h11 == _t_T_34[15:8] ? 8'h82 : _GEN_4112; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4114 = 8'h12 == _t_T_34[15:8] ? 8'hc9 : _GEN_4113; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4115 = 8'h13 == _t_T_34[15:8] ? 8'h7d : _GEN_4114; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4116 = 8'h14 == _t_T_34[15:8] ? 8'hfa : _GEN_4115; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4117 = 8'h15 == _t_T_34[15:8] ? 8'h59 : _GEN_4116; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4118 = 8'h16 == _t_T_34[15:8] ? 8'h47 : _GEN_4117; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4119 = 8'h17 == _t_T_34[15:8] ? 8'hf0 : _GEN_4118; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4120 = 8'h18 == _t_T_34[15:8] ? 8'had : _GEN_4119; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4121 = 8'h19 == _t_T_34[15:8] ? 8'hd4 : _GEN_4120; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4122 = 8'h1a == _t_T_34[15:8] ? 8'ha2 : _GEN_4121; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4123 = 8'h1b == _t_T_34[15:8] ? 8'haf : _GEN_4122; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4124 = 8'h1c == _t_T_34[15:8] ? 8'h9c : _GEN_4123; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4125 = 8'h1d == _t_T_34[15:8] ? 8'ha4 : _GEN_4124; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4126 = 8'h1e == _t_T_34[15:8] ? 8'h72 : _GEN_4125; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4127 = 8'h1f == _t_T_34[15:8] ? 8'hc0 : _GEN_4126; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4128 = 8'h20 == _t_T_34[15:8] ? 8'hb7 : _GEN_4127; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4129 = 8'h21 == _t_T_34[15:8] ? 8'hfd : _GEN_4128; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4130 = 8'h22 == _t_T_34[15:8] ? 8'h93 : _GEN_4129; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4131 = 8'h23 == _t_T_34[15:8] ? 8'h26 : _GEN_4130; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4132 = 8'h24 == _t_T_34[15:8] ? 8'h36 : _GEN_4131; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4133 = 8'h25 == _t_T_34[15:8] ? 8'h3f : _GEN_4132; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4134 = 8'h26 == _t_T_34[15:8] ? 8'hf7 : _GEN_4133; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4135 = 8'h27 == _t_T_34[15:8] ? 8'hcc : _GEN_4134; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4136 = 8'h28 == _t_T_34[15:8] ? 8'h34 : _GEN_4135; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4137 = 8'h29 == _t_T_34[15:8] ? 8'ha5 : _GEN_4136; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4138 = 8'h2a == _t_T_34[15:8] ? 8'he5 : _GEN_4137; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4139 = 8'h2b == _t_T_34[15:8] ? 8'hf1 : _GEN_4138; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4140 = 8'h2c == _t_T_34[15:8] ? 8'h71 : _GEN_4139; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4141 = 8'h2d == _t_T_34[15:8] ? 8'hd8 : _GEN_4140; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4142 = 8'h2e == _t_T_34[15:8] ? 8'h31 : _GEN_4141; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4143 = 8'h2f == _t_T_34[15:8] ? 8'h15 : _GEN_4142; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4144 = 8'h30 == _t_T_34[15:8] ? 8'h4 : _GEN_4143; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4145 = 8'h31 == _t_T_34[15:8] ? 8'hc7 : _GEN_4144; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4146 = 8'h32 == _t_T_34[15:8] ? 8'h23 : _GEN_4145; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4147 = 8'h33 == _t_T_34[15:8] ? 8'hc3 : _GEN_4146; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4148 = 8'h34 == _t_T_34[15:8] ? 8'h18 : _GEN_4147; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4149 = 8'h35 == _t_T_34[15:8] ? 8'h96 : _GEN_4148; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4150 = 8'h36 == _t_T_34[15:8] ? 8'h5 : _GEN_4149; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4151 = 8'h37 == _t_T_34[15:8] ? 8'h9a : _GEN_4150; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4152 = 8'h38 == _t_T_34[15:8] ? 8'h7 : _GEN_4151; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4153 = 8'h39 == _t_T_34[15:8] ? 8'h12 : _GEN_4152; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4154 = 8'h3a == _t_T_34[15:8] ? 8'h80 : _GEN_4153; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4155 = 8'h3b == _t_T_34[15:8] ? 8'he2 : _GEN_4154; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4156 = 8'h3c == _t_T_34[15:8] ? 8'heb : _GEN_4155; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4157 = 8'h3d == _t_T_34[15:8] ? 8'h27 : _GEN_4156; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4158 = 8'h3e == _t_T_34[15:8] ? 8'hb2 : _GEN_4157; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4159 = 8'h3f == _t_T_34[15:8] ? 8'h75 : _GEN_4158; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4160 = 8'h40 == _t_T_34[15:8] ? 8'h9 : _GEN_4159; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4161 = 8'h41 == _t_T_34[15:8] ? 8'h83 : _GEN_4160; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4162 = 8'h42 == _t_T_34[15:8] ? 8'h2c : _GEN_4161; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4163 = 8'h43 == _t_T_34[15:8] ? 8'h1a : _GEN_4162; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4164 = 8'h44 == _t_T_34[15:8] ? 8'h1b : _GEN_4163; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4165 = 8'h45 == _t_T_34[15:8] ? 8'h6e : _GEN_4164; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4166 = 8'h46 == _t_T_34[15:8] ? 8'h5a : _GEN_4165; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4167 = 8'h47 == _t_T_34[15:8] ? 8'ha0 : _GEN_4166; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4168 = 8'h48 == _t_T_34[15:8] ? 8'h52 : _GEN_4167; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4169 = 8'h49 == _t_T_34[15:8] ? 8'h3b : _GEN_4168; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4170 = 8'h4a == _t_T_34[15:8] ? 8'hd6 : _GEN_4169; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4171 = 8'h4b == _t_T_34[15:8] ? 8'hb3 : _GEN_4170; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4172 = 8'h4c == _t_T_34[15:8] ? 8'h29 : _GEN_4171; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4173 = 8'h4d == _t_T_34[15:8] ? 8'he3 : _GEN_4172; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4174 = 8'h4e == _t_T_34[15:8] ? 8'h2f : _GEN_4173; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4175 = 8'h4f == _t_T_34[15:8] ? 8'h84 : _GEN_4174; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4176 = 8'h50 == _t_T_34[15:8] ? 8'h53 : _GEN_4175; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4177 = 8'h51 == _t_T_34[15:8] ? 8'hd1 : _GEN_4176; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4178 = 8'h52 == _t_T_34[15:8] ? 8'h0 : _GEN_4177; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4179 = 8'h53 == _t_T_34[15:8] ? 8'hed : _GEN_4178; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4180 = 8'h54 == _t_T_34[15:8] ? 8'h20 : _GEN_4179; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4181 = 8'h55 == _t_T_34[15:8] ? 8'hfc : _GEN_4180; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4182 = 8'h56 == _t_T_34[15:8] ? 8'hb1 : _GEN_4181; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4183 = 8'h57 == _t_T_34[15:8] ? 8'h5b : _GEN_4182; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4184 = 8'h58 == _t_T_34[15:8] ? 8'h6a : _GEN_4183; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4185 = 8'h59 == _t_T_34[15:8] ? 8'hcb : _GEN_4184; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4186 = 8'h5a == _t_T_34[15:8] ? 8'hbe : _GEN_4185; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4187 = 8'h5b == _t_T_34[15:8] ? 8'h39 : _GEN_4186; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4188 = 8'h5c == _t_T_34[15:8] ? 8'h4a : _GEN_4187; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4189 = 8'h5d == _t_T_34[15:8] ? 8'h4c : _GEN_4188; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4190 = 8'h5e == _t_T_34[15:8] ? 8'h58 : _GEN_4189; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4191 = 8'h5f == _t_T_34[15:8] ? 8'hcf : _GEN_4190; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4192 = 8'h60 == _t_T_34[15:8] ? 8'hd0 : _GEN_4191; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4193 = 8'h61 == _t_T_34[15:8] ? 8'hef : _GEN_4192; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4194 = 8'h62 == _t_T_34[15:8] ? 8'haa : _GEN_4193; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4195 = 8'h63 == _t_T_34[15:8] ? 8'hfb : _GEN_4194; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4196 = 8'h64 == _t_T_34[15:8] ? 8'h43 : _GEN_4195; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4197 = 8'h65 == _t_T_34[15:8] ? 8'h4d : _GEN_4196; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4198 = 8'h66 == _t_T_34[15:8] ? 8'h33 : _GEN_4197; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4199 = 8'h67 == _t_T_34[15:8] ? 8'h85 : _GEN_4198; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4200 = 8'h68 == _t_T_34[15:8] ? 8'h45 : _GEN_4199; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4201 = 8'h69 == _t_T_34[15:8] ? 8'hf9 : _GEN_4200; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4202 = 8'h6a == _t_T_34[15:8] ? 8'h2 : _GEN_4201; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4203 = 8'h6b == _t_T_34[15:8] ? 8'h7f : _GEN_4202; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4204 = 8'h6c == _t_T_34[15:8] ? 8'h50 : _GEN_4203; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4205 = 8'h6d == _t_T_34[15:8] ? 8'h3c : _GEN_4204; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4206 = 8'h6e == _t_T_34[15:8] ? 8'h9f : _GEN_4205; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4207 = 8'h6f == _t_T_34[15:8] ? 8'ha8 : _GEN_4206; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4208 = 8'h70 == _t_T_34[15:8] ? 8'h51 : _GEN_4207; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4209 = 8'h71 == _t_T_34[15:8] ? 8'ha3 : _GEN_4208; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4210 = 8'h72 == _t_T_34[15:8] ? 8'h40 : _GEN_4209; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4211 = 8'h73 == _t_T_34[15:8] ? 8'h8f : _GEN_4210; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4212 = 8'h74 == _t_T_34[15:8] ? 8'h92 : _GEN_4211; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4213 = 8'h75 == _t_T_34[15:8] ? 8'h9d : _GEN_4212; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4214 = 8'h76 == _t_T_34[15:8] ? 8'h38 : _GEN_4213; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4215 = 8'h77 == _t_T_34[15:8] ? 8'hf5 : _GEN_4214; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4216 = 8'h78 == _t_T_34[15:8] ? 8'hbc : _GEN_4215; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4217 = 8'h79 == _t_T_34[15:8] ? 8'hb6 : _GEN_4216; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4218 = 8'h7a == _t_T_34[15:8] ? 8'hda : _GEN_4217; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4219 = 8'h7b == _t_T_34[15:8] ? 8'h21 : _GEN_4218; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4220 = 8'h7c == _t_T_34[15:8] ? 8'h10 : _GEN_4219; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4221 = 8'h7d == _t_T_34[15:8] ? 8'hff : _GEN_4220; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4222 = 8'h7e == _t_T_34[15:8] ? 8'hf3 : _GEN_4221; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4223 = 8'h7f == _t_T_34[15:8] ? 8'hd2 : _GEN_4222; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4224 = 8'h80 == _t_T_34[15:8] ? 8'hcd : _GEN_4223; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4225 = 8'h81 == _t_T_34[15:8] ? 8'hc : _GEN_4224; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4226 = 8'h82 == _t_T_34[15:8] ? 8'h13 : _GEN_4225; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4227 = 8'h83 == _t_T_34[15:8] ? 8'hec : _GEN_4226; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4228 = 8'h84 == _t_T_34[15:8] ? 8'h5f : _GEN_4227; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4229 = 8'h85 == _t_T_34[15:8] ? 8'h97 : _GEN_4228; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4230 = 8'h86 == _t_T_34[15:8] ? 8'h44 : _GEN_4229; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4231 = 8'h87 == _t_T_34[15:8] ? 8'h17 : _GEN_4230; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4232 = 8'h88 == _t_T_34[15:8] ? 8'hc4 : _GEN_4231; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4233 = 8'h89 == _t_T_34[15:8] ? 8'ha7 : _GEN_4232; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4234 = 8'h8a == _t_T_34[15:8] ? 8'h7e : _GEN_4233; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4235 = 8'h8b == _t_T_34[15:8] ? 8'h3d : _GEN_4234; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4236 = 8'h8c == _t_T_34[15:8] ? 8'h64 : _GEN_4235; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4237 = 8'h8d == _t_T_34[15:8] ? 8'h5d : _GEN_4236; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4238 = 8'h8e == _t_T_34[15:8] ? 8'h19 : _GEN_4237; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4239 = 8'h8f == _t_T_34[15:8] ? 8'h73 : _GEN_4238; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4240 = 8'h90 == _t_T_34[15:8] ? 8'h60 : _GEN_4239; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4241 = 8'h91 == _t_T_34[15:8] ? 8'h81 : _GEN_4240; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4242 = 8'h92 == _t_T_34[15:8] ? 8'h4f : _GEN_4241; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4243 = 8'h93 == _t_T_34[15:8] ? 8'hdc : _GEN_4242; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4244 = 8'h94 == _t_T_34[15:8] ? 8'h22 : _GEN_4243; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4245 = 8'h95 == _t_T_34[15:8] ? 8'h2a : _GEN_4244; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4246 = 8'h96 == _t_T_34[15:8] ? 8'h90 : _GEN_4245; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4247 = 8'h97 == _t_T_34[15:8] ? 8'h88 : _GEN_4246; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4248 = 8'h98 == _t_T_34[15:8] ? 8'h46 : _GEN_4247; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4249 = 8'h99 == _t_T_34[15:8] ? 8'hee : _GEN_4248; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4250 = 8'h9a == _t_T_34[15:8] ? 8'hb8 : _GEN_4249; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4251 = 8'h9b == _t_T_34[15:8] ? 8'h14 : _GEN_4250; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4252 = 8'h9c == _t_T_34[15:8] ? 8'hde : _GEN_4251; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4253 = 8'h9d == _t_T_34[15:8] ? 8'h5e : _GEN_4252; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4254 = 8'h9e == _t_T_34[15:8] ? 8'hb : _GEN_4253; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4255 = 8'h9f == _t_T_34[15:8] ? 8'hdb : _GEN_4254; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4256 = 8'ha0 == _t_T_34[15:8] ? 8'he0 : _GEN_4255; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4257 = 8'ha1 == _t_T_34[15:8] ? 8'h32 : _GEN_4256; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4258 = 8'ha2 == _t_T_34[15:8] ? 8'h3a : _GEN_4257; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4259 = 8'ha3 == _t_T_34[15:8] ? 8'ha : _GEN_4258; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4260 = 8'ha4 == _t_T_34[15:8] ? 8'h49 : _GEN_4259; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4261 = 8'ha5 == _t_T_34[15:8] ? 8'h6 : _GEN_4260; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4262 = 8'ha6 == _t_T_34[15:8] ? 8'h24 : _GEN_4261; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4263 = 8'ha7 == _t_T_34[15:8] ? 8'h5c : _GEN_4262; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4264 = 8'ha8 == _t_T_34[15:8] ? 8'hc2 : _GEN_4263; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4265 = 8'ha9 == _t_T_34[15:8] ? 8'hd3 : _GEN_4264; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4266 = 8'haa == _t_T_34[15:8] ? 8'hac : _GEN_4265; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4267 = 8'hab == _t_T_34[15:8] ? 8'h62 : _GEN_4266; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4268 = 8'hac == _t_T_34[15:8] ? 8'h91 : _GEN_4267; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4269 = 8'had == _t_T_34[15:8] ? 8'h95 : _GEN_4268; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4270 = 8'hae == _t_T_34[15:8] ? 8'he4 : _GEN_4269; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4271 = 8'haf == _t_T_34[15:8] ? 8'h79 : _GEN_4270; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4272 = 8'hb0 == _t_T_34[15:8] ? 8'he7 : _GEN_4271; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4273 = 8'hb1 == _t_T_34[15:8] ? 8'hc8 : _GEN_4272; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4274 = 8'hb2 == _t_T_34[15:8] ? 8'h37 : _GEN_4273; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4275 = 8'hb3 == _t_T_34[15:8] ? 8'h6d : _GEN_4274; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4276 = 8'hb4 == _t_T_34[15:8] ? 8'h8d : _GEN_4275; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4277 = 8'hb5 == _t_T_34[15:8] ? 8'hd5 : _GEN_4276; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4278 = 8'hb6 == _t_T_34[15:8] ? 8'h4e : _GEN_4277; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4279 = 8'hb7 == _t_T_34[15:8] ? 8'ha9 : _GEN_4278; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4280 = 8'hb8 == _t_T_34[15:8] ? 8'h6c : _GEN_4279; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4281 = 8'hb9 == _t_T_34[15:8] ? 8'h56 : _GEN_4280; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4282 = 8'hba == _t_T_34[15:8] ? 8'hf4 : _GEN_4281; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4283 = 8'hbb == _t_T_34[15:8] ? 8'hea : _GEN_4282; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4284 = 8'hbc == _t_T_34[15:8] ? 8'h65 : _GEN_4283; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4285 = 8'hbd == _t_T_34[15:8] ? 8'h7a : _GEN_4284; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4286 = 8'hbe == _t_T_34[15:8] ? 8'hae : _GEN_4285; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4287 = 8'hbf == _t_T_34[15:8] ? 8'h8 : _GEN_4286; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4288 = 8'hc0 == _t_T_34[15:8] ? 8'hba : _GEN_4287; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4289 = 8'hc1 == _t_T_34[15:8] ? 8'h78 : _GEN_4288; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4290 = 8'hc2 == _t_T_34[15:8] ? 8'h25 : _GEN_4289; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4291 = 8'hc3 == _t_T_34[15:8] ? 8'h2e : _GEN_4290; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4292 = 8'hc4 == _t_T_34[15:8] ? 8'h1c : _GEN_4291; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4293 = 8'hc5 == _t_T_34[15:8] ? 8'ha6 : _GEN_4292; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4294 = 8'hc6 == _t_T_34[15:8] ? 8'hb4 : _GEN_4293; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4295 = 8'hc7 == _t_T_34[15:8] ? 8'hc6 : _GEN_4294; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4296 = 8'hc8 == _t_T_34[15:8] ? 8'he8 : _GEN_4295; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4297 = 8'hc9 == _t_T_34[15:8] ? 8'hdd : _GEN_4296; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4298 = 8'hca == _t_T_34[15:8] ? 8'h74 : _GEN_4297; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4299 = 8'hcb == _t_T_34[15:8] ? 8'h1f : _GEN_4298; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4300 = 8'hcc == _t_T_34[15:8] ? 8'h4b : _GEN_4299; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4301 = 8'hcd == _t_T_34[15:8] ? 8'hbd : _GEN_4300; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4302 = 8'hce == _t_T_34[15:8] ? 8'h8b : _GEN_4301; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4303 = 8'hcf == _t_T_34[15:8] ? 8'h8a : _GEN_4302; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4304 = 8'hd0 == _t_T_34[15:8] ? 8'h70 : _GEN_4303; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4305 = 8'hd1 == _t_T_34[15:8] ? 8'h3e : _GEN_4304; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4306 = 8'hd2 == _t_T_34[15:8] ? 8'hb5 : _GEN_4305; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4307 = 8'hd3 == _t_T_34[15:8] ? 8'h66 : _GEN_4306; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4308 = 8'hd4 == _t_T_34[15:8] ? 8'h48 : _GEN_4307; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4309 = 8'hd5 == _t_T_34[15:8] ? 8'h3 : _GEN_4308; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4310 = 8'hd6 == _t_T_34[15:8] ? 8'hf6 : _GEN_4309; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4311 = 8'hd7 == _t_T_34[15:8] ? 8'he : _GEN_4310; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4312 = 8'hd8 == _t_T_34[15:8] ? 8'h61 : _GEN_4311; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4313 = 8'hd9 == _t_T_34[15:8] ? 8'h35 : _GEN_4312; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4314 = 8'hda == _t_T_34[15:8] ? 8'h57 : _GEN_4313; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4315 = 8'hdb == _t_T_34[15:8] ? 8'hb9 : _GEN_4314; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4316 = 8'hdc == _t_T_34[15:8] ? 8'h86 : _GEN_4315; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4317 = 8'hdd == _t_T_34[15:8] ? 8'hc1 : _GEN_4316; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4318 = 8'hde == _t_T_34[15:8] ? 8'h1d : _GEN_4317; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4319 = 8'hdf == _t_T_34[15:8] ? 8'h9e : _GEN_4318; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4320 = 8'he0 == _t_T_34[15:8] ? 8'he1 : _GEN_4319; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4321 = 8'he1 == _t_T_34[15:8] ? 8'hf8 : _GEN_4320; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4322 = 8'he2 == _t_T_34[15:8] ? 8'h98 : _GEN_4321; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4323 = 8'he3 == _t_T_34[15:8] ? 8'h11 : _GEN_4322; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4324 = 8'he4 == _t_T_34[15:8] ? 8'h69 : _GEN_4323; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4325 = 8'he5 == _t_T_34[15:8] ? 8'hd9 : _GEN_4324; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4326 = 8'he6 == _t_T_34[15:8] ? 8'h8e : _GEN_4325; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4327 = 8'he7 == _t_T_34[15:8] ? 8'h94 : _GEN_4326; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4328 = 8'he8 == _t_T_34[15:8] ? 8'h9b : _GEN_4327; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4329 = 8'he9 == _t_T_34[15:8] ? 8'h1e : _GEN_4328; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4330 = 8'hea == _t_T_34[15:8] ? 8'h87 : _GEN_4329; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4331 = 8'heb == _t_T_34[15:8] ? 8'he9 : _GEN_4330; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4332 = 8'hec == _t_T_34[15:8] ? 8'hce : _GEN_4331; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4333 = 8'hed == _t_T_34[15:8] ? 8'h55 : _GEN_4332; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4334 = 8'hee == _t_T_34[15:8] ? 8'h28 : _GEN_4333; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4335 = 8'hef == _t_T_34[15:8] ? 8'hdf : _GEN_4334; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4336 = 8'hf0 == _t_T_34[15:8] ? 8'h8c : _GEN_4335; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4337 = 8'hf1 == _t_T_34[15:8] ? 8'ha1 : _GEN_4336; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4338 = 8'hf2 == _t_T_34[15:8] ? 8'h89 : _GEN_4337; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4339 = 8'hf3 == _t_T_34[15:8] ? 8'hd : _GEN_4338; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4340 = 8'hf4 == _t_T_34[15:8] ? 8'hbf : _GEN_4339; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4341 = 8'hf5 == _t_T_34[15:8] ? 8'he6 : _GEN_4340; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4342 = 8'hf6 == _t_T_34[15:8] ? 8'h42 : _GEN_4341; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4343 = 8'hf7 == _t_T_34[15:8] ? 8'h68 : _GEN_4342; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4344 = 8'hf8 == _t_T_34[15:8] ? 8'h41 : _GEN_4343; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4345 = 8'hf9 == _t_T_34[15:8] ? 8'h99 : _GEN_4344; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4346 = 8'hfa == _t_T_34[15:8] ? 8'h2d : _GEN_4345; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4347 = 8'hfb == _t_T_34[15:8] ? 8'hf : _GEN_4346; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4348 = 8'hfc == _t_T_34[15:8] ? 8'hb0 : _GEN_4347; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4349 = 8'hfd == _t_T_34[15:8] ? 8'h54 : _GEN_4348; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4350 = 8'hfe == _t_T_34[15:8] ? 8'hbb : _GEN_4349; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4351 = 8'hff == _t_T_34[15:8] ? 8'h16 : _GEN_4350; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4353 = 8'h1 == _t_T_34[7:0] ? 8'h7c : 8'h63; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4354 = 8'h2 == _t_T_34[7:0] ? 8'h77 : _GEN_4353; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4355 = 8'h3 == _t_T_34[7:0] ? 8'h7b : _GEN_4354; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4356 = 8'h4 == _t_T_34[7:0] ? 8'hf2 : _GEN_4355; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4357 = 8'h5 == _t_T_34[7:0] ? 8'h6b : _GEN_4356; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4358 = 8'h6 == _t_T_34[7:0] ? 8'h6f : _GEN_4357; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4359 = 8'h7 == _t_T_34[7:0] ? 8'hc5 : _GEN_4358; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4360 = 8'h8 == _t_T_34[7:0] ? 8'h30 : _GEN_4359; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4361 = 8'h9 == _t_T_34[7:0] ? 8'h1 : _GEN_4360; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4362 = 8'ha == _t_T_34[7:0] ? 8'h67 : _GEN_4361; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4363 = 8'hb == _t_T_34[7:0] ? 8'h2b : _GEN_4362; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4364 = 8'hc == _t_T_34[7:0] ? 8'hfe : _GEN_4363; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4365 = 8'hd == _t_T_34[7:0] ? 8'hd7 : _GEN_4364; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4366 = 8'he == _t_T_34[7:0] ? 8'hab : _GEN_4365; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4367 = 8'hf == _t_T_34[7:0] ? 8'h76 : _GEN_4366; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4368 = 8'h10 == _t_T_34[7:0] ? 8'hca : _GEN_4367; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4369 = 8'h11 == _t_T_34[7:0] ? 8'h82 : _GEN_4368; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4370 = 8'h12 == _t_T_34[7:0] ? 8'hc9 : _GEN_4369; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4371 = 8'h13 == _t_T_34[7:0] ? 8'h7d : _GEN_4370; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4372 = 8'h14 == _t_T_34[7:0] ? 8'hfa : _GEN_4371; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4373 = 8'h15 == _t_T_34[7:0] ? 8'h59 : _GEN_4372; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4374 = 8'h16 == _t_T_34[7:0] ? 8'h47 : _GEN_4373; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4375 = 8'h17 == _t_T_34[7:0] ? 8'hf0 : _GEN_4374; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4376 = 8'h18 == _t_T_34[7:0] ? 8'had : _GEN_4375; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4377 = 8'h19 == _t_T_34[7:0] ? 8'hd4 : _GEN_4376; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4378 = 8'h1a == _t_T_34[7:0] ? 8'ha2 : _GEN_4377; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4379 = 8'h1b == _t_T_34[7:0] ? 8'haf : _GEN_4378; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4380 = 8'h1c == _t_T_34[7:0] ? 8'h9c : _GEN_4379; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4381 = 8'h1d == _t_T_34[7:0] ? 8'ha4 : _GEN_4380; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4382 = 8'h1e == _t_T_34[7:0] ? 8'h72 : _GEN_4381; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4383 = 8'h1f == _t_T_34[7:0] ? 8'hc0 : _GEN_4382; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4384 = 8'h20 == _t_T_34[7:0] ? 8'hb7 : _GEN_4383; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4385 = 8'h21 == _t_T_34[7:0] ? 8'hfd : _GEN_4384; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4386 = 8'h22 == _t_T_34[7:0] ? 8'h93 : _GEN_4385; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4387 = 8'h23 == _t_T_34[7:0] ? 8'h26 : _GEN_4386; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4388 = 8'h24 == _t_T_34[7:0] ? 8'h36 : _GEN_4387; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4389 = 8'h25 == _t_T_34[7:0] ? 8'h3f : _GEN_4388; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4390 = 8'h26 == _t_T_34[7:0] ? 8'hf7 : _GEN_4389; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4391 = 8'h27 == _t_T_34[7:0] ? 8'hcc : _GEN_4390; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4392 = 8'h28 == _t_T_34[7:0] ? 8'h34 : _GEN_4391; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4393 = 8'h29 == _t_T_34[7:0] ? 8'ha5 : _GEN_4392; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4394 = 8'h2a == _t_T_34[7:0] ? 8'he5 : _GEN_4393; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4395 = 8'h2b == _t_T_34[7:0] ? 8'hf1 : _GEN_4394; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4396 = 8'h2c == _t_T_34[7:0] ? 8'h71 : _GEN_4395; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4397 = 8'h2d == _t_T_34[7:0] ? 8'hd8 : _GEN_4396; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4398 = 8'h2e == _t_T_34[7:0] ? 8'h31 : _GEN_4397; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4399 = 8'h2f == _t_T_34[7:0] ? 8'h15 : _GEN_4398; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4400 = 8'h30 == _t_T_34[7:0] ? 8'h4 : _GEN_4399; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4401 = 8'h31 == _t_T_34[7:0] ? 8'hc7 : _GEN_4400; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4402 = 8'h32 == _t_T_34[7:0] ? 8'h23 : _GEN_4401; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4403 = 8'h33 == _t_T_34[7:0] ? 8'hc3 : _GEN_4402; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4404 = 8'h34 == _t_T_34[7:0] ? 8'h18 : _GEN_4403; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4405 = 8'h35 == _t_T_34[7:0] ? 8'h96 : _GEN_4404; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4406 = 8'h36 == _t_T_34[7:0] ? 8'h5 : _GEN_4405; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4407 = 8'h37 == _t_T_34[7:0] ? 8'h9a : _GEN_4406; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4408 = 8'h38 == _t_T_34[7:0] ? 8'h7 : _GEN_4407; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4409 = 8'h39 == _t_T_34[7:0] ? 8'h12 : _GEN_4408; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4410 = 8'h3a == _t_T_34[7:0] ? 8'h80 : _GEN_4409; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4411 = 8'h3b == _t_T_34[7:0] ? 8'he2 : _GEN_4410; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4412 = 8'h3c == _t_T_34[7:0] ? 8'heb : _GEN_4411; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4413 = 8'h3d == _t_T_34[7:0] ? 8'h27 : _GEN_4412; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4414 = 8'h3e == _t_T_34[7:0] ? 8'hb2 : _GEN_4413; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4415 = 8'h3f == _t_T_34[7:0] ? 8'h75 : _GEN_4414; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4416 = 8'h40 == _t_T_34[7:0] ? 8'h9 : _GEN_4415; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4417 = 8'h41 == _t_T_34[7:0] ? 8'h83 : _GEN_4416; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4418 = 8'h42 == _t_T_34[7:0] ? 8'h2c : _GEN_4417; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4419 = 8'h43 == _t_T_34[7:0] ? 8'h1a : _GEN_4418; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4420 = 8'h44 == _t_T_34[7:0] ? 8'h1b : _GEN_4419; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4421 = 8'h45 == _t_T_34[7:0] ? 8'h6e : _GEN_4420; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4422 = 8'h46 == _t_T_34[7:0] ? 8'h5a : _GEN_4421; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4423 = 8'h47 == _t_T_34[7:0] ? 8'ha0 : _GEN_4422; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4424 = 8'h48 == _t_T_34[7:0] ? 8'h52 : _GEN_4423; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4425 = 8'h49 == _t_T_34[7:0] ? 8'h3b : _GEN_4424; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4426 = 8'h4a == _t_T_34[7:0] ? 8'hd6 : _GEN_4425; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4427 = 8'h4b == _t_T_34[7:0] ? 8'hb3 : _GEN_4426; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4428 = 8'h4c == _t_T_34[7:0] ? 8'h29 : _GEN_4427; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4429 = 8'h4d == _t_T_34[7:0] ? 8'he3 : _GEN_4428; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4430 = 8'h4e == _t_T_34[7:0] ? 8'h2f : _GEN_4429; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4431 = 8'h4f == _t_T_34[7:0] ? 8'h84 : _GEN_4430; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4432 = 8'h50 == _t_T_34[7:0] ? 8'h53 : _GEN_4431; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4433 = 8'h51 == _t_T_34[7:0] ? 8'hd1 : _GEN_4432; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4434 = 8'h52 == _t_T_34[7:0] ? 8'h0 : _GEN_4433; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4435 = 8'h53 == _t_T_34[7:0] ? 8'hed : _GEN_4434; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4436 = 8'h54 == _t_T_34[7:0] ? 8'h20 : _GEN_4435; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4437 = 8'h55 == _t_T_34[7:0] ? 8'hfc : _GEN_4436; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4438 = 8'h56 == _t_T_34[7:0] ? 8'hb1 : _GEN_4437; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4439 = 8'h57 == _t_T_34[7:0] ? 8'h5b : _GEN_4438; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4440 = 8'h58 == _t_T_34[7:0] ? 8'h6a : _GEN_4439; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4441 = 8'h59 == _t_T_34[7:0] ? 8'hcb : _GEN_4440; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4442 = 8'h5a == _t_T_34[7:0] ? 8'hbe : _GEN_4441; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4443 = 8'h5b == _t_T_34[7:0] ? 8'h39 : _GEN_4442; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4444 = 8'h5c == _t_T_34[7:0] ? 8'h4a : _GEN_4443; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4445 = 8'h5d == _t_T_34[7:0] ? 8'h4c : _GEN_4444; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4446 = 8'h5e == _t_T_34[7:0] ? 8'h58 : _GEN_4445; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4447 = 8'h5f == _t_T_34[7:0] ? 8'hcf : _GEN_4446; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4448 = 8'h60 == _t_T_34[7:0] ? 8'hd0 : _GEN_4447; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4449 = 8'h61 == _t_T_34[7:0] ? 8'hef : _GEN_4448; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4450 = 8'h62 == _t_T_34[7:0] ? 8'haa : _GEN_4449; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4451 = 8'h63 == _t_T_34[7:0] ? 8'hfb : _GEN_4450; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4452 = 8'h64 == _t_T_34[7:0] ? 8'h43 : _GEN_4451; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4453 = 8'h65 == _t_T_34[7:0] ? 8'h4d : _GEN_4452; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4454 = 8'h66 == _t_T_34[7:0] ? 8'h33 : _GEN_4453; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4455 = 8'h67 == _t_T_34[7:0] ? 8'h85 : _GEN_4454; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4456 = 8'h68 == _t_T_34[7:0] ? 8'h45 : _GEN_4455; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4457 = 8'h69 == _t_T_34[7:0] ? 8'hf9 : _GEN_4456; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4458 = 8'h6a == _t_T_34[7:0] ? 8'h2 : _GEN_4457; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4459 = 8'h6b == _t_T_34[7:0] ? 8'h7f : _GEN_4458; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4460 = 8'h6c == _t_T_34[7:0] ? 8'h50 : _GEN_4459; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4461 = 8'h6d == _t_T_34[7:0] ? 8'h3c : _GEN_4460; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4462 = 8'h6e == _t_T_34[7:0] ? 8'h9f : _GEN_4461; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4463 = 8'h6f == _t_T_34[7:0] ? 8'ha8 : _GEN_4462; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4464 = 8'h70 == _t_T_34[7:0] ? 8'h51 : _GEN_4463; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4465 = 8'h71 == _t_T_34[7:0] ? 8'ha3 : _GEN_4464; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4466 = 8'h72 == _t_T_34[7:0] ? 8'h40 : _GEN_4465; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4467 = 8'h73 == _t_T_34[7:0] ? 8'h8f : _GEN_4466; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4468 = 8'h74 == _t_T_34[7:0] ? 8'h92 : _GEN_4467; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4469 = 8'h75 == _t_T_34[7:0] ? 8'h9d : _GEN_4468; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4470 = 8'h76 == _t_T_34[7:0] ? 8'h38 : _GEN_4469; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4471 = 8'h77 == _t_T_34[7:0] ? 8'hf5 : _GEN_4470; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4472 = 8'h78 == _t_T_34[7:0] ? 8'hbc : _GEN_4471; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4473 = 8'h79 == _t_T_34[7:0] ? 8'hb6 : _GEN_4472; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4474 = 8'h7a == _t_T_34[7:0] ? 8'hda : _GEN_4473; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4475 = 8'h7b == _t_T_34[7:0] ? 8'h21 : _GEN_4474; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4476 = 8'h7c == _t_T_34[7:0] ? 8'h10 : _GEN_4475; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4477 = 8'h7d == _t_T_34[7:0] ? 8'hff : _GEN_4476; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4478 = 8'h7e == _t_T_34[7:0] ? 8'hf3 : _GEN_4477; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4479 = 8'h7f == _t_T_34[7:0] ? 8'hd2 : _GEN_4478; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4480 = 8'h80 == _t_T_34[7:0] ? 8'hcd : _GEN_4479; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4481 = 8'h81 == _t_T_34[7:0] ? 8'hc : _GEN_4480; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4482 = 8'h82 == _t_T_34[7:0] ? 8'h13 : _GEN_4481; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4483 = 8'h83 == _t_T_34[7:0] ? 8'hec : _GEN_4482; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4484 = 8'h84 == _t_T_34[7:0] ? 8'h5f : _GEN_4483; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4485 = 8'h85 == _t_T_34[7:0] ? 8'h97 : _GEN_4484; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4486 = 8'h86 == _t_T_34[7:0] ? 8'h44 : _GEN_4485; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4487 = 8'h87 == _t_T_34[7:0] ? 8'h17 : _GEN_4486; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4488 = 8'h88 == _t_T_34[7:0] ? 8'hc4 : _GEN_4487; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4489 = 8'h89 == _t_T_34[7:0] ? 8'ha7 : _GEN_4488; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4490 = 8'h8a == _t_T_34[7:0] ? 8'h7e : _GEN_4489; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4491 = 8'h8b == _t_T_34[7:0] ? 8'h3d : _GEN_4490; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4492 = 8'h8c == _t_T_34[7:0] ? 8'h64 : _GEN_4491; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4493 = 8'h8d == _t_T_34[7:0] ? 8'h5d : _GEN_4492; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4494 = 8'h8e == _t_T_34[7:0] ? 8'h19 : _GEN_4493; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4495 = 8'h8f == _t_T_34[7:0] ? 8'h73 : _GEN_4494; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4496 = 8'h90 == _t_T_34[7:0] ? 8'h60 : _GEN_4495; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4497 = 8'h91 == _t_T_34[7:0] ? 8'h81 : _GEN_4496; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4498 = 8'h92 == _t_T_34[7:0] ? 8'h4f : _GEN_4497; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4499 = 8'h93 == _t_T_34[7:0] ? 8'hdc : _GEN_4498; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4500 = 8'h94 == _t_T_34[7:0] ? 8'h22 : _GEN_4499; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4501 = 8'h95 == _t_T_34[7:0] ? 8'h2a : _GEN_4500; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4502 = 8'h96 == _t_T_34[7:0] ? 8'h90 : _GEN_4501; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4503 = 8'h97 == _t_T_34[7:0] ? 8'h88 : _GEN_4502; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4504 = 8'h98 == _t_T_34[7:0] ? 8'h46 : _GEN_4503; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4505 = 8'h99 == _t_T_34[7:0] ? 8'hee : _GEN_4504; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4506 = 8'h9a == _t_T_34[7:0] ? 8'hb8 : _GEN_4505; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4507 = 8'h9b == _t_T_34[7:0] ? 8'h14 : _GEN_4506; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4508 = 8'h9c == _t_T_34[7:0] ? 8'hde : _GEN_4507; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4509 = 8'h9d == _t_T_34[7:0] ? 8'h5e : _GEN_4508; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4510 = 8'h9e == _t_T_34[7:0] ? 8'hb : _GEN_4509; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4511 = 8'h9f == _t_T_34[7:0] ? 8'hdb : _GEN_4510; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4512 = 8'ha0 == _t_T_34[7:0] ? 8'he0 : _GEN_4511; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4513 = 8'ha1 == _t_T_34[7:0] ? 8'h32 : _GEN_4512; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4514 = 8'ha2 == _t_T_34[7:0] ? 8'h3a : _GEN_4513; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4515 = 8'ha3 == _t_T_34[7:0] ? 8'ha : _GEN_4514; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4516 = 8'ha4 == _t_T_34[7:0] ? 8'h49 : _GEN_4515; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4517 = 8'ha5 == _t_T_34[7:0] ? 8'h6 : _GEN_4516; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4518 = 8'ha6 == _t_T_34[7:0] ? 8'h24 : _GEN_4517; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4519 = 8'ha7 == _t_T_34[7:0] ? 8'h5c : _GEN_4518; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4520 = 8'ha8 == _t_T_34[7:0] ? 8'hc2 : _GEN_4519; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4521 = 8'ha9 == _t_T_34[7:0] ? 8'hd3 : _GEN_4520; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4522 = 8'haa == _t_T_34[7:0] ? 8'hac : _GEN_4521; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4523 = 8'hab == _t_T_34[7:0] ? 8'h62 : _GEN_4522; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4524 = 8'hac == _t_T_34[7:0] ? 8'h91 : _GEN_4523; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4525 = 8'had == _t_T_34[7:0] ? 8'h95 : _GEN_4524; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4526 = 8'hae == _t_T_34[7:0] ? 8'he4 : _GEN_4525; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4527 = 8'haf == _t_T_34[7:0] ? 8'h79 : _GEN_4526; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4528 = 8'hb0 == _t_T_34[7:0] ? 8'he7 : _GEN_4527; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4529 = 8'hb1 == _t_T_34[7:0] ? 8'hc8 : _GEN_4528; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4530 = 8'hb2 == _t_T_34[7:0] ? 8'h37 : _GEN_4529; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4531 = 8'hb3 == _t_T_34[7:0] ? 8'h6d : _GEN_4530; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4532 = 8'hb4 == _t_T_34[7:0] ? 8'h8d : _GEN_4531; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4533 = 8'hb5 == _t_T_34[7:0] ? 8'hd5 : _GEN_4532; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4534 = 8'hb6 == _t_T_34[7:0] ? 8'h4e : _GEN_4533; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4535 = 8'hb7 == _t_T_34[7:0] ? 8'ha9 : _GEN_4534; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4536 = 8'hb8 == _t_T_34[7:0] ? 8'h6c : _GEN_4535; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4537 = 8'hb9 == _t_T_34[7:0] ? 8'h56 : _GEN_4536; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4538 = 8'hba == _t_T_34[7:0] ? 8'hf4 : _GEN_4537; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4539 = 8'hbb == _t_T_34[7:0] ? 8'hea : _GEN_4538; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4540 = 8'hbc == _t_T_34[7:0] ? 8'h65 : _GEN_4539; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4541 = 8'hbd == _t_T_34[7:0] ? 8'h7a : _GEN_4540; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4542 = 8'hbe == _t_T_34[7:0] ? 8'hae : _GEN_4541; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4543 = 8'hbf == _t_T_34[7:0] ? 8'h8 : _GEN_4542; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4544 = 8'hc0 == _t_T_34[7:0] ? 8'hba : _GEN_4543; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4545 = 8'hc1 == _t_T_34[7:0] ? 8'h78 : _GEN_4544; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4546 = 8'hc2 == _t_T_34[7:0] ? 8'h25 : _GEN_4545; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4547 = 8'hc3 == _t_T_34[7:0] ? 8'h2e : _GEN_4546; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4548 = 8'hc4 == _t_T_34[7:0] ? 8'h1c : _GEN_4547; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4549 = 8'hc5 == _t_T_34[7:0] ? 8'ha6 : _GEN_4548; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4550 = 8'hc6 == _t_T_34[7:0] ? 8'hb4 : _GEN_4549; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4551 = 8'hc7 == _t_T_34[7:0] ? 8'hc6 : _GEN_4550; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4552 = 8'hc8 == _t_T_34[7:0] ? 8'he8 : _GEN_4551; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4553 = 8'hc9 == _t_T_34[7:0] ? 8'hdd : _GEN_4552; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4554 = 8'hca == _t_T_34[7:0] ? 8'h74 : _GEN_4553; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4555 = 8'hcb == _t_T_34[7:0] ? 8'h1f : _GEN_4554; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4556 = 8'hcc == _t_T_34[7:0] ? 8'h4b : _GEN_4555; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4557 = 8'hcd == _t_T_34[7:0] ? 8'hbd : _GEN_4556; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4558 = 8'hce == _t_T_34[7:0] ? 8'h8b : _GEN_4557; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4559 = 8'hcf == _t_T_34[7:0] ? 8'h8a : _GEN_4558; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4560 = 8'hd0 == _t_T_34[7:0] ? 8'h70 : _GEN_4559; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4561 = 8'hd1 == _t_T_34[7:0] ? 8'h3e : _GEN_4560; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4562 = 8'hd2 == _t_T_34[7:0] ? 8'hb5 : _GEN_4561; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4563 = 8'hd3 == _t_T_34[7:0] ? 8'h66 : _GEN_4562; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4564 = 8'hd4 == _t_T_34[7:0] ? 8'h48 : _GEN_4563; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4565 = 8'hd5 == _t_T_34[7:0] ? 8'h3 : _GEN_4564; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4566 = 8'hd6 == _t_T_34[7:0] ? 8'hf6 : _GEN_4565; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4567 = 8'hd7 == _t_T_34[7:0] ? 8'he : _GEN_4566; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4568 = 8'hd8 == _t_T_34[7:0] ? 8'h61 : _GEN_4567; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4569 = 8'hd9 == _t_T_34[7:0] ? 8'h35 : _GEN_4568; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4570 = 8'hda == _t_T_34[7:0] ? 8'h57 : _GEN_4569; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4571 = 8'hdb == _t_T_34[7:0] ? 8'hb9 : _GEN_4570; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4572 = 8'hdc == _t_T_34[7:0] ? 8'h86 : _GEN_4571; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4573 = 8'hdd == _t_T_34[7:0] ? 8'hc1 : _GEN_4572; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4574 = 8'hde == _t_T_34[7:0] ? 8'h1d : _GEN_4573; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4575 = 8'hdf == _t_T_34[7:0] ? 8'h9e : _GEN_4574; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4576 = 8'he0 == _t_T_34[7:0] ? 8'he1 : _GEN_4575; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4577 = 8'he1 == _t_T_34[7:0] ? 8'hf8 : _GEN_4576; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4578 = 8'he2 == _t_T_34[7:0] ? 8'h98 : _GEN_4577; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4579 = 8'he3 == _t_T_34[7:0] ? 8'h11 : _GEN_4578; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4580 = 8'he4 == _t_T_34[7:0] ? 8'h69 : _GEN_4579; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4581 = 8'he5 == _t_T_34[7:0] ? 8'hd9 : _GEN_4580; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4582 = 8'he6 == _t_T_34[7:0] ? 8'h8e : _GEN_4581; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4583 = 8'he7 == _t_T_34[7:0] ? 8'h94 : _GEN_4582; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4584 = 8'he8 == _t_T_34[7:0] ? 8'h9b : _GEN_4583; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4585 = 8'he9 == _t_T_34[7:0] ? 8'h1e : _GEN_4584; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4586 = 8'hea == _t_T_34[7:0] ? 8'h87 : _GEN_4585; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4587 = 8'heb == _t_T_34[7:0] ? 8'he9 : _GEN_4586; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4588 = 8'hec == _t_T_34[7:0] ? 8'hce : _GEN_4587; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4589 = 8'hed == _t_T_34[7:0] ? 8'h55 : _GEN_4588; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4590 = 8'hee == _t_T_34[7:0] ? 8'h28 : _GEN_4589; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4591 = 8'hef == _t_T_34[7:0] ? 8'hdf : _GEN_4590; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4592 = 8'hf0 == _t_T_34[7:0] ? 8'h8c : _GEN_4591; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4593 = 8'hf1 == _t_T_34[7:0] ? 8'ha1 : _GEN_4592; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4594 = 8'hf2 == _t_T_34[7:0] ? 8'h89 : _GEN_4593; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4595 = 8'hf3 == _t_T_34[7:0] ? 8'hd : _GEN_4594; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4596 = 8'hf4 == _t_T_34[7:0] ? 8'hbf : _GEN_4595; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4597 = 8'hf5 == _t_T_34[7:0] ? 8'he6 : _GEN_4596; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4598 = 8'hf6 == _t_T_34[7:0] ? 8'h42 : _GEN_4597; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4599 = 8'hf7 == _t_T_34[7:0] ? 8'h68 : _GEN_4598; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4600 = 8'hf8 == _t_T_34[7:0] ? 8'h41 : _GEN_4599; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4601 = 8'hf9 == _t_T_34[7:0] ? 8'h99 : _GEN_4600; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4602 = 8'hfa == _t_T_34[7:0] ? 8'h2d : _GEN_4601; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4603 = 8'hfb == _t_T_34[7:0] ? 8'hf : _GEN_4602; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4604 = 8'hfc == _t_T_34[7:0] ? 8'hb0 : _GEN_4603; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4605 = 8'hfd == _t_T_34[7:0] ? 8'h54 : _GEN_4604; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4606 = 8'hfe == _t_T_34[7:0] ? 8'hbb : _GEN_4605; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4607 = 8'hff == _t_T_34[7:0] ? 8'h16 : _GEN_4606; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4609 = 8'h1 == _t_T_34[31:24] ? 8'h7c : 8'h63; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4610 = 8'h2 == _t_T_34[31:24] ? 8'h77 : _GEN_4609; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4611 = 8'h3 == _t_T_34[31:24] ? 8'h7b : _GEN_4610; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4612 = 8'h4 == _t_T_34[31:24] ? 8'hf2 : _GEN_4611; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4613 = 8'h5 == _t_T_34[31:24] ? 8'h6b : _GEN_4612; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4614 = 8'h6 == _t_T_34[31:24] ? 8'h6f : _GEN_4613; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4615 = 8'h7 == _t_T_34[31:24] ? 8'hc5 : _GEN_4614; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4616 = 8'h8 == _t_T_34[31:24] ? 8'h30 : _GEN_4615; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4617 = 8'h9 == _t_T_34[31:24] ? 8'h1 : _GEN_4616; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4618 = 8'ha == _t_T_34[31:24] ? 8'h67 : _GEN_4617; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4619 = 8'hb == _t_T_34[31:24] ? 8'h2b : _GEN_4618; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4620 = 8'hc == _t_T_34[31:24] ? 8'hfe : _GEN_4619; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4621 = 8'hd == _t_T_34[31:24] ? 8'hd7 : _GEN_4620; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4622 = 8'he == _t_T_34[31:24] ? 8'hab : _GEN_4621; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4623 = 8'hf == _t_T_34[31:24] ? 8'h76 : _GEN_4622; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4624 = 8'h10 == _t_T_34[31:24] ? 8'hca : _GEN_4623; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4625 = 8'h11 == _t_T_34[31:24] ? 8'h82 : _GEN_4624; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4626 = 8'h12 == _t_T_34[31:24] ? 8'hc9 : _GEN_4625; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4627 = 8'h13 == _t_T_34[31:24] ? 8'h7d : _GEN_4626; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4628 = 8'h14 == _t_T_34[31:24] ? 8'hfa : _GEN_4627; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4629 = 8'h15 == _t_T_34[31:24] ? 8'h59 : _GEN_4628; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4630 = 8'h16 == _t_T_34[31:24] ? 8'h47 : _GEN_4629; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4631 = 8'h17 == _t_T_34[31:24] ? 8'hf0 : _GEN_4630; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4632 = 8'h18 == _t_T_34[31:24] ? 8'had : _GEN_4631; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4633 = 8'h19 == _t_T_34[31:24] ? 8'hd4 : _GEN_4632; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4634 = 8'h1a == _t_T_34[31:24] ? 8'ha2 : _GEN_4633; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4635 = 8'h1b == _t_T_34[31:24] ? 8'haf : _GEN_4634; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4636 = 8'h1c == _t_T_34[31:24] ? 8'h9c : _GEN_4635; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4637 = 8'h1d == _t_T_34[31:24] ? 8'ha4 : _GEN_4636; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4638 = 8'h1e == _t_T_34[31:24] ? 8'h72 : _GEN_4637; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4639 = 8'h1f == _t_T_34[31:24] ? 8'hc0 : _GEN_4638; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4640 = 8'h20 == _t_T_34[31:24] ? 8'hb7 : _GEN_4639; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4641 = 8'h21 == _t_T_34[31:24] ? 8'hfd : _GEN_4640; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4642 = 8'h22 == _t_T_34[31:24] ? 8'h93 : _GEN_4641; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4643 = 8'h23 == _t_T_34[31:24] ? 8'h26 : _GEN_4642; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4644 = 8'h24 == _t_T_34[31:24] ? 8'h36 : _GEN_4643; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4645 = 8'h25 == _t_T_34[31:24] ? 8'h3f : _GEN_4644; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4646 = 8'h26 == _t_T_34[31:24] ? 8'hf7 : _GEN_4645; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4647 = 8'h27 == _t_T_34[31:24] ? 8'hcc : _GEN_4646; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4648 = 8'h28 == _t_T_34[31:24] ? 8'h34 : _GEN_4647; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4649 = 8'h29 == _t_T_34[31:24] ? 8'ha5 : _GEN_4648; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4650 = 8'h2a == _t_T_34[31:24] ? 8'he5 : _GEN_4649; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4651 = 8'h2b == _t_T_34[31:24] ? 8'hf1 : _GEN_4650; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4652 = 8'h2c == _t_T_34[31:24] ? 8'h71 : _GEN_4651; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4653 = 8'h2d == _t_T_34[31:24] ? 8'hd8 : _GEN_4652; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4654 = 8'h2e == _t_T_34[31:24] ? 8'h31 : _GEN_4653; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4655 = 8'h2f == _t_T_34[31:24] ? 8'h15 : _GEN_4654; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4656 = 8'h30 == _t_T_34[31:24] ? 8'h4 : _GEN_4655; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4657 = 8'h31 == _t_T_34[31:24] ? 8'hc7 : _GEN_4656; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4658 = 8'h32 == _t_T_34[31:24] ? 8'h23 : _GEN_4657; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4659 = 8'h33 == _t_T_34[31:24] ? 8'hc3 : _GEN_4658; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4660 = 8'h34 == _t_T_34[31:24] ? 8'h18 : _GEN_4659; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4661 = 8'h35 == _t_T_34[31:24] ? 8'h96 : _GEN_4660; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4662 = 8'h36 == _t_T_34[31:24] ? 8'h5 : _GEN_4661; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4663 = 8'h37 == _t_T_34[31:24] ? 8'h9a : _GEN_4662; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4664 = 8'h38 == _t_T_34[31:24] ? 8'h7 : _GEN_4663; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4665 = 8'h39 == _t_T_34[31:24] ? 8'h12 : _GEN_4664; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4666 = 8'h3a == _t_T_34[31:24] ? 8'h80 : _GEN_4665; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4667 = 8'h3b == _t_T_34[31:24] ? 8'he2 : _GEN_4666; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4668 = 8'h3c == _t_T_34[31:24] ? 8'heb : _GEN_4667; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4669 = 8'h3d == _t_T_34[31:24] ? 8'h27 : _GEN_4668; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4670 = 8'h3e == _t_T_34[31:24] ? 8'hb2 : _GEN_4669; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4671 = 8'h3f == _t_T_34[31:24] ? 8'h75 : _GEN_4670; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4672 = 8'h40 == _t_T_34[31:24] ? 8'h9 : _GEN_4671; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4673 = 8'h41 == _t_T_34[31:24] ? 8'h83 : _GEN_4672; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4674 = 8'h42 == _t_T_34[31:24] ? 8'h2c : _GEN_4673; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4675 = 8'h43 == _t_T_34[31:24] ? 8'h1a : _GEN_4674; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4676 = 8'h44 == _t_T_34[31:24] ? 8'h1b : _GEN_4675; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4677 = 8'h45 == _t_T_34[31:24] ? 8'h6e : _GEN_4676; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4678 = 8'h46 == _t_T_34[31:24] ? 8'h5a : _GEN_4677; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4679 = 8'h47 == _t_T_34[31:24] ? 8'ha0 : _GEN_4678; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4680 = 8'h48 == _t_T_34[31:24] ? 8'h52 : _GEN_4679; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4681 = 8'h49 == _t_T_34[31:24] ? 8'h3b : _GEN_4680; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4682 = 8'h4a == _t_T_34[31:24] ? 8'hd6 : _GEN_4681; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4683 = 8'h4b == _t_T_34[31:24] ? 8'hb3 : _GEN_4682; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4684 = 8'h4c == _t_T_34[31:24] ? 8'h29 : _GEN_4683; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4685 = 8'h4d == _t_T_34[31:24] ? 8'he3 : _GEN_4684; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4686 = 8'h4e == _t_T_34[31:24] ? 8'h2f : _GEN_4685; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4687 = 8'h4f == _t_T_34[31:24] ? 8'h84 : _GEN_4686; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4688 = 8'h50 == _t_T_34[31:24] ? 8'h53 : _GEN_4687; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4689 = 8'h51 == _t_T_34[31:24] ? 8'hd1 : _GEN_4688; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4690 = 8'h52 == _t_T_34[31:24] ? 8'h0 : _GEN_4689; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4691 = 8'h53 == _t_T_34[31:24] ? 8'hed : _GEN_4690; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4692 = 8'h54 == _t_T_34[31:24] ? 8'h20 : _GEN_4691; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4693 = 8'h55 == _t_T_34[31:24] ? 8'hfc : _GEN_4692; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4694 = 8'h56 == _t_T_34[31:24] ? 8'hb1 : _GEN_4693; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4695 = 8'h57 == _t_T_34[31:24] ? 8'h5b : _GEN_4694; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4696 = 8'h58 == _t_T_34[31:24] ? 8'h6a : _GEN_4695; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4697 = 8'h59 == _t_T_34[31:24] ? 8'hcb : _GEN_4696; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4698 = 8'h5a == _t_T_34[31:24] ? 8'hbe : _GEN_4697; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4699 = 8'h5b == _t_T_34[31:24] ? 8'h39 : _GEN_4698; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4700 = 8'h5c == _t_T_34[31:24] ? 8'h4a : _GEN_4699; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4701 = 8'h5d == _t_T_34[31:24] ? 8'h4c : _GEN_4700; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4702 = 8'h5e == _t_T_34[31:24] ? 8'h58 : _GEN_4701; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4703 = 8'h5f == _t_T_34[31:24] ? 8'hcf : _GEN_4702; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4704 = 8'h60 == _t_T_34[31:24] ? 8'hd0 : _GEN_4703; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4705 = 8'h61 == _t_T_34[31:24] ? 8'hef : _GEN_4704; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4706 = 8'h62 == _t_T_34[31:24] ? 8'haa : _GEN_4705; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4707 = 8'h63 == _t_T_34[31:24] ? 8'hfb : _GEN_4706; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4708 = 8'h64 == _t_T_34[31:24] ? 8'h43 : _GEN_4707; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4709 = 8'h65 == _t_T_34[31:24] ? 8'h4d : _GEN_4708; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4710 = 8'h66 == _t_T_34[31:24] ? 8'h33 : _GEN_4709; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4711 = 8'h67 == _t_T_34[31:24] ? 8'h85 : _GEN_4710; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4712 = 8'h68 == _t_T_34[31:24] ? 8'h45 : _GEN_4711; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4713 = 8'h69 == _t_T_34[31:24] ? 8'hf9 : _GEN_4712; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4714 = 8'h6a == _t_T_34[31:24] ? 8'h2 : _GEN_4713; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4715 = 8'h6b == _t_T_34[31:24] ? 8'h7f : _GEN_4714; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4716 = 8'h6c == _t_T_34[31:24] ? 8'h50 : _GEN_4715; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4717 = 8'h6d == _t_T_34[31:24] ? 8'h3c : _GEN_4716; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4718 = 8'h6e == _t_T_34[31:24] ? 8'h9f : _GEN_4717; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4719 = 8'h6f == _t_T_34[31:24] ? 8'ha8 : _GEN_4718; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4720 = 8'h70 == _t_T_34[31:24] ? 8'h51 : _GEN_4719; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4721 = 8'h71 == _t_T_34[31:24] ? 8'ha3 : _GEN_4720; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4722 = 8'h72 == _t_T_34[31:24] ? 8'h40 : _GEN_4721; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4723 = 8'h73 == _t_T_34[31:24] ? 8'h8f : _GEN_4722; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4724 = 8'h74 == _t_T_34[31:24] ? 8'h92 : _GEN_4723; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4725 = 8'h75 == _t_T_34[31:24] ? 8'h9d : _GEN_4724; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4726 = 8'h76 == _t_T_34[31:24] ? 8'h38 : _GEN_4725; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4727 = 8'h77 == _t_T_34[31:24] ? 8'hf5 : _GEN_4726; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4728 = 8'h78 == _t_T_34[31:24] ? 8'hbc : _GEN_4727; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4729 = 8'h79 == _t_T_34[31:24] ? 8'hb6 : _GEN_4728; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4730 = 8'h7a == _t_T_34[31:24] ? 8'hda : _GEN_4729; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4731 = 8'h7b == _t_T_34[31:24] ? 8'h21 : _GEN_4730; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4732 = 8'h7c == _t_T_34[31:24] ? 8'h10 : _GEN_4731; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4733 = 8'h7d == _t_T_34[31:24] ? 8'hff : _GEN_4732; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4734 = 8'h7e == _t_T_34[31:24] ? 8'hf3 : _GEN_4733; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4735 = 8'h7f == _t_T_34[31:24] ? 8'hd2 : _GEN_4734; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4736 = 8'h80 == _t_T_34[31:24] ? 8'hcd : _GEN_4735; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4737 = 8'h81 == _t_T_34[31:24] ? 8'hc : _GEN_4736; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4738 = 8'h82 == _t_T_34[31:24] ? 8'h13 : _GEN_4737; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4739 = 8'h83 == _t_T_34[31:24] ? 8'hec : _GEN_4738; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4740 = 8'h84 == _t_T_34[31:24] ? 8'h5f : _GEN_4739; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4741 = 8'h85 == _t_T_34[31:24] ? 8'h97 : _GEN_4740; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4742 = 8'h86 == _t_T_34[31:24] ? 8'h44 : _GEN_4741; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4743 = 8'h87 == _t_T_34[31:24] ? 8'h17 : _GEN_4742; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4744 = 8'h88 == _t_T_34[31:24] ? 8'hc4 : _GEN_4743; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4745 = 8'h89 == _t_T_34[31:24] ? 8'ha7 : _GEN_4744; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4746 = 8'h8a == _t_T_34[31:24] ? 8'h7e : _GEN_4745; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4747 = 8'h8b == _t_T_34[31:24] ? 8'h3d : _GEN_4746; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4748 = 8'h8c == _t_T_34[31:24] ? 8'h64 : _GEN_4747; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4749 = 8'h8d == _t_T_34[31:24] ? 8'h5d : _GEN_4748; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4750 = 8'h8e == _t_T_34[31:24] ? 8'h19 : _GEN_4749; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4751 = 8'h8f == _t_T_34[31:24] ? 8'h73 : _GEN_4750; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4752 = 8'h90 == _t_T_34[31:24] ? 8'h60 : _GEN_4751; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4753 = 8'h91 == _t_T_34[31:24] ? 8'h81 : _GEN_4752; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4754 = 8'h92 == _t_T_34[31:24] ? 8'h4f : _GEN_4753; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4755 = 8'h93 == _t_T_34[31:24] ? 8'hdc : _GEN_4754; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4756 = 8'h94 == _t_T_34[31:24] ? 8'h22 : _GEN_4755; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4757 = 8'h95 == _t_T_34[31:24] ? 8'h2a : _GEN_4756; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4758 = 8'h96 == _t_T_34[31:24] ? 8'h90 : _GEN_4757; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4759 = 8'h97 == _t_T_34[31:24] ? 8'h88 : _GEN_4758; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4760 = 8'h98 == _t_T_34[31:24] ? 8'h46 : _GEN_4759; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4761 = 8'h99 == _t_T_34[31:24] ? 8'hee : _GEN_4760; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4762 = 8'h9a == _t_T_34[31:24] ? 8'hb8 : _GEN_4761; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4763 = 8'h9b == _t_T_34[31:24] ? 8'h14 : _GEN_4762; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4764 = 8'h9c == _t_T_34[31:24] ? 8'hde : _GEN_4763; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4765 = 8'h9d == _t_T_34[31:24] ? 8'h5e : _GEN_4764; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4766 = 8'h9e == _t_T_34[31:24] ? 8'hb : _GEN_4765; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4767 = 8'h9f == _t_T_34[31:24] ? 8'hdb : _GEN_4766; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4768 = 8'ha0 == _t_T_34[31:24] ? 8'he0 : _GEN_4767; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4769 = 8'ha1 == _t_T_34[31:24] ? 8'h32 : _GEN_4768; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4770 = 8'ha2 == _t_T_34[31:24] ? 8'h3a : _GEN_4769; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4771 = 8'ha3 == _t_T_34[31:24] ? 8'ha : _GEN_4770; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4772 = 8'ha4 == _t_T_34[31:24] ? 8'h49 : _GEN_4771; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4773 = 8'ha5 == _t_T_34[31:24] ? 8'h6 : _GEN_4772; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4774 = 8'ha6 == _t_T_34[31:24] ? 8'h24 : _GEN_4773; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4775 = 8'ha7 == _t_T_34[31:24] ? 8'h5c : _GEN_4774; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4776 = 8'ha8 == _t_T_34[31:24] ? 8'hc2 : _GEN_4775; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4777 = 8'ha9 == _t_T_34[31:24] ? 8'hd3 : _GEN_4776; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4778 = 8'haa == _t_T_34[31:24] ? 8'hac : _GEN_4777; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4779 = 8'hab == _t_T_34[31:24] ? 8'h62 : _GEN_4778; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4780 = 8'hac == _t_T_34[31:24] ? 8'h91 : _GEN_4779; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4781 = 8'had == _t_T_34[31:24] ? 8'h95 : _GEN_4780; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4782 = 8'hae == _t_T_34[31:24] ? 8'he4 : _GEN_4781; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4783 = 8'haf == _t_T_34[31:24] ? 8'h79 : _GEN_4782; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4784 = 8'hb0 == _t_T_34[31:24] ? 8'he7 : _GEN_4783; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4785 = 8'hb1 == _t_T_34[31:24] ? 8'hc8 : _GEN_4784; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4786 = 8'hb2 == _t_T_34[31:24] ? 8'h37 : _GEN_4785; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4787 = 8'hb3 == _t_T_34[31:24] ? 8'h6d : _GEN_4786; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4788 = 8'hb4 == _t_T_34[31:24] ? 8'h8d : _GEN_4787; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4789 = 8'hb5 == _t_T_34[31:24] ? 8'hd5 : _GEN_4788; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4790 = 8'hb6 == _t_T_34[31:24] ? 8'h4e : _GEN_4789; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4791 = 8'hb7 == _t_T_34[31:24] ? 8'ha9 : _GEN_4790; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4792 = 8'hb8 == _t_T_34[31:24] ? 8'h6c : _GEN_4791; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4793 = 8'hb9 == _t_T_34[31:24] ? 8'h56 : _GEN_4792; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4794 = 8'hba == _t_T_34[31:24] ? 8'hf4 : _GEN_4793; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4795 = 8'hbb == _t_T_34[31:24] ? 8'hea : _GEN_4794; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4796 = 8'hbc == _t_T_34[31:24] ? 8'h65 : _GEN_4795; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4797 = 8'hbd == _t_T_34[31:24] ? 8'h7a : _GEN_4796; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4798 = 8'hbe == _t_T_34[31:24] ? 8'hae : _GEN_4797; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4799 = 8'hbf == _t_T_34[31:24] ? 8'h8 : _GEN_4798; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4800 = 8'hc0 == _t_T_34[31:24] ? 8'hba : _GEN_4799; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4801 = 8'hc1 == _t_T_34[31:24] ? 8'h78 : _GEN_4800; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4802 = 8'hc2 == _t_T_34[31:24] ? 8'h25 : _GEN_4801; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4803 = 8'hc3 == _t_T_34[31:24] ? 8'h2e : _GEN_4802; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4804 = 8'hc4 == _t_T_34[31:24] ? 8'h1c : _GEN_4803; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4805 = 8'hc5 == _t_T_34[31:24] ? 8'ha6 : _GEN_4804; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4806 = 8'hc6 == _t_T_34[31:24] ? 8'hb4 : _GEN_4805; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4807 = 8'hc7 == _t_T_34[31:24] ? 8'hc6 : _GEN_4806; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4808 = 8'hc8 == _t_T_34[31:24] ? 8'he8 : _GEN_4807; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4809 = 8'hc9 == _t_T_34[31:24] ? 8'hdd : _GEN_4808; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4810 = 8'hca == _t_T_34[31:24] ? 8'h74 : _GEN_4809; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4811 = 8'hcb == _t_T_34[31:24] ? 8'h1f : _GEN_4810; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4812 = 8'hcc == _t_T_34[31:24] ? 8'h4b : _GEN_4811; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4813 = 8'hcd == _t_T_34[31:24] ? 8'hbd : _GEN_4812; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4814 = 8'hce == _t_T_34[31:24] ? 8'h8b : _GEN_4813; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4815 = 8'hcf == _t_T_34[31:24] ? 8'h8a : _GEN_4814; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4816 = 8'hd0 == _t_T_34[31:24] ? 8'h70 : _GEN_4815; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4817 = 8'hd1 == _t_T_34[31:24] ? 8'h3e : _GEN_4816; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4818 = 8'hd2 == _t_T_34[31:24] ? 8'hb5 : _GEN_4817; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4819 = 8'hd3 == _t_T_34[31:24] ? 8'h66 : _GEN_4818; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4820 = 8'hd4 == _t_T_34[31:24] ? 8'h48 : _GEN_4819; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4821 = 8'hd5 == _t_T_34[31:24] ? 8'h3 : _GEN_4820; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4822 = 8'hd6 == _t_T_34[31:24] ? 8'hf6 : _GEN_4821; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4823 = 8'hd7 == _t_T_34[31:24] ? 8'he : _GEN_4822; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4824 = 8'hd8 == _t_T_34[31:24] ? 8'h61 : _GEN_4823; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4825 = 8'hd9 == _t_T_34[31:24] ? 8'h35 : _GEN_4824; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4826 = 8'hda == _t_T_34[31:24] ? 8'h57 : _GEN_4825; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4827 = 8'hdb == _t_T_34[31:24] ? 8'hb9 : _GEN_4826; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4828 = 8'hdc == _t_T_34[31:24] ? 8'h86 : _GEN_4827; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4829 = 8'hdd == _t_T_34[31:24] ? 8'hc1 : _GEN_4828; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4830 = 8'hde == _t_T_34[31:24] ? 8'h1d : _GEN_4829; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4831 = 8'hdf == _t_T_34[31:24] ? 8'h9e : _GEN_4830; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4832 = 8'he0 == _t_T_34[31:24] ? 8'he1 : _GEN_4831; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4833 = 8'he1 == _t_T_34[31:24] ? 8'hf8 : _GEN_4832; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4834 = 8'he2 == _t_T_34[31:24] ? 8'h98 : _GEN_4833; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4835 = 8'he3 == _t_T_34[31:24] ? 8'h11 : _GEN_4834; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4836 = 8'he4 == _t_T_34[31:24] ? 8'h69 : _GEN_4835; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4837 = 8'he5 == _t_T_34[31:24] ? 8'hd9 : _GEN_4836; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4838 = 8'he6 == _t_T_34[31:24] ? 8'h8e : _GEN_4837; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4839 = 8'he7 == _t_T_34[31:24] ? 8'h94 : _GEN_4838; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4840 = 8'he8 == _t_T_34[31:24] ? 8'h9b : _GEN_4839; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4841 = 8'he9 == _t_T_34[31:24] ? 8'h1e : _GEN_4840; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4842 = 8'hea == _t_T_34[31:24] ? 8'h87 : _GEN_4841; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4843 = 8'heb == _t_T_34[31:24] ? 8'he9 : _GEN_4842; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4844 = 8'hec == _t_T_34[31:24] ? 8'hce : _GEN_4843; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4845 = 8'hed == _t_T_34[31:24] ? 8'h55 : _GEN_4844; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4846 = 8'hee == _t_T_34[31:24] ? 8'h28 : _GEN_4845; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4847 = 8'hef == _t_T_34[31:24] ? 8'hdf : _GEN_4846; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4848 = 8'hf0 == _t_T_34[31:24] ? 8'h8c : _GEN_4847; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4849 = 8'hf1 == _t_T_34[31:24] ? 8'ha1 : _GEN_4848; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4850 = 8'hf2 == _t_T_34[31:24] ? 8'h89 : _GEN_4849; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4851 = 8'hf3 == _t_T_34[31:24] ? 8'hd : _GEN_4850; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4852 = 8'hf4 == _t_T_34[31:24] ? 8'hbf : _GEN_4851; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4853 = 8'hf5 == _t_T_34[31:24] ? 8'he6 : _GEN_4852; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4854 = 8'hf6 == _t_T_34[31:24] ? 8'h42 : _GEN_4853; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4855 = 8'hf7 == _t_T_34[31:24] ? 8'h68 : _GEN_4854; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4856 = 8'hf8 == _t_T_34[31:24] ? 8'h41 : _GEN_4855; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4857 = 8'hf9 == _t_T_34[31:24] ? 8'h99 : _GEN_4856; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4858 = 8'hfa == _t_T_34[31:24] ? 8'h2d : _GEN_4857; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4859 = 8'hfb == _t_T_34[31:24] ? 8'hf : _GEN_4858; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4860 = 8'hfc == _t_T_34[31:24] ? 8'hb0 : _GEN_4859; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4861 = 8'hfd == _t_T_34[31:24] ? 8'h54 : _GEN_4860; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4862 = 8'hfe == _t_T_34[31:24] ? 8'hbb : _GEN_4861; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4863 = 8'hff == _t_T_34[31:24] ? 8'h16 : _GEN_4862; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4865 = 8'h1 == _t_T_34[23:16] ? 8'h7c : 8'h63; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4866 = 8'h2 == _t_T_34[23:16] ? 8'h77 : _GEN_4865; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4867 = 8'h3 == _t_T_34[23:16] ? 8'h7b : _GEN_4866; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4868 = 8'h4 == _t_T_34[23:16] ? 8'hf2 : _GEN_4867; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4869 = 8'h5 == _t_T_34[23:16] ? 8'h6b : _GEN_4868; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4870 = 8'h6 == _t_T_34[23:16] ? 8'h6f : _GEN_4869; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4871 = 8'h7 == _t_T_34[23:16] ? 8'hc5 : _GEN_4870; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4872 = 8'h8 == _t_T_34[23:16] ? 8'h30 : _GEN_4871; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4873 = 8'h9 == _t_T_34[23:16] ? 8'h1 : _GEN_4872; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4874 = 8'ha == _t_T_34[23:16] ? 8'h67 : _GEN_4873; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4875 = 8'hb == _t_T_34[23:16] ? 8'h2b : _GEN_4874; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4876 = 8'hc == _t_T_34[23:16] ? 8'hfe : _GEN_4875; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4877 = 8'hd == _t_T_34[23:16] ? 8'hd7 : _GEN_4876; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4878 = 8'he == _t_T_34[23:16] ? 8'hab : _GEN_4877; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4879 = 8'hf == _t_T_34[23:16] ? 8'h76 : _GEN_4878; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4880 = 8'h10 == _t_T_34[23:16] ? 8'hca : _GEN_4879; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4881 = 8'h11 == _t_T_34[23:16] ? 8'h82 : _GEN_4880; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4882 = 8'h12 == _t_T_34[23:16] ? 8'hc9 : _GEN_4881; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4883 = 8'h13 == _t_T_34[23:16] ? 8'h7d : _GEN_4882; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4884 = 8'h14 == _t_T_34[23:16] ? 8'hfa : _GEN_4883; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4885 = 8'h15 == _t_T_34[23:16] ? 8'h59 : _GEN_4884; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4886 = 8'h16 == _t_T_34[23:16] ? 8'h47 : _GEN_4885; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4887 = 8'h17 == _t_T_34[23:16] ? 8'hf0 : _GEN_4886; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4888 = 8'h18 == _t_T_34[23:16] ? 8'had : _GEN_4887; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4889 = 8'h19 == _t_T_34[23:16] ? 8'hd4 : _GEN_4888; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4890 = 8'h1a == _t_T_34[23:16] ? 8'ha2 : _GEN_4889; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4891 = 8'h1b == _t_T_34[23:16] ? 8'haf : _GEN_4890; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4892 = 8'h1c == _t_T_34[23:16] ? 8'h9c : _GEN_4891; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4893 = 8'h1d == _t_T_34[23:16] ? 8'ha4 : _GEN_4892; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4894 = 8'h1e == _t_T_34[23:16] ? 8'h72 : _GEN_4893; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4895 = 8'h1f == _t_T_34[23:16] ? 8'hc0 : _GEN_4894; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4896 = 8'h20 == _t_T_34[23:16] ? 8'hb7 : _GEN_4895; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4897 = 8'h21 == _t_T_34[23:16] ? 8'hfd : _GEN_4896; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4898 = 8'h22 == _t_T_34[23:16] ? 8'h93 : _GEN_4897; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4899 = 8'h23 == _t_T_34[23:16] ? 8'h26 : _GEN_4898; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4900 = 8'h24 == _t_T_34[23:16] ? 8'h36 : _GEN_4899; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4901 = 8'h25 == _t_T_34[23:16] ? 8'h3f : _GEN_4900; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4902 = 8'h26 == _t_T_34[23:16] ? 8'hf7 : _GEN_4901; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4903 = 8'h27 == _t_T_34[23:16] ? 8'hcc : _GEN_4902; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4904 = 8'h28 == _t_T_34[23:16] ? 8'h34 : _GEN_4903; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4905 = 8'h29 == _t_T_34[23:16] ? 8'ha5 : _GEN_4904; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4906 = 8'h2a == _t_T_34[23:16] ? 8'he5 : _GEN_4905; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4907 = 8'h2b == _t_T_34[23:16] ? 8'hf1 : _GEN_4906; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4908 = 8'h2c == _t_T_34[23:16] ? 8'h71 : _GEN_4907; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4909 = 8'h2d == _t_T_34[23:16] ? 8'hd8 : _GEN_4908; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4910 = 8'h2e == _t_T_34[23:16] ? 8'h31 : _GEN_4909; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4911 = 8'h2f == _t_T_34[23:16] ? 8'h15 : _GEN_4910; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4912 = 8'h30 == _t_T_34[23:16] ? 8'h4 : _GEN_4911; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4913 = 8'h31 == _t_T_34[23:16] ? 8'hc7 : _GEN_4912; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4914 = 8'h32 == _t_T_34[23:16] ? 8'h23 : _GEN_4913; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4915 = 8'h33 == _t_T_34[23:16] ? 8'hc3 : _GEN_4914; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4916 = 8'h34 == _t_T_34[23:16] ? 8'h18 : _GEN_4915; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4917 = 8'h35 == _t_T_34[23:16] ? 8'h96 : _GEN_4916; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4918 = 8'h36 == _t_T_34[23:16] ? 8'h5 : _GEN_4917; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4919 = 8'h37 == _t_T_34[23:16] ? 8'h9a : _GEN_4918; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4920 = 8'h38 == _t_T_34[23:16] ? 8'h7 : _GEN_4919; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4921 = 8'h39 == _t_T_34[23:16] ? 8'h12 : _GEN_4920; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4922 = 8'h3a == _t_T_34[23:16] ? 8'h80 : _GEN_4921; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4923 = 8'h3b == _t_T_34[23:16] ? 8'he2 : _GEN_4922; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4924 = 8'h3c == _t_T_34[23:16] ? 8'heb : _GEN_4923; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4925 = 8'h3d == _t_T_34[23:16] ? 8'h27 : _GEN_4924; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4926 = 8'h3e == _t_T_34[23:16] ? 8'hb2 : _GEN_4925; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4927 = 8'h3f == _t_T_34[23:16] ? 8'h75 : _GEN_4926; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4928 = 8'h40 == _t_T_34[23:16] ? 8'h9 : _GEN_4927; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4929 = 8'h41 == _t_T_34[23:16] ? 8'h83 : _GEN_4928; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4930 = 8'h42 == _t_T_34[23:16] ? 8'h2c : _GEN_4929; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4931 = 8'h43 == _t_T_34[23:16] ? 8'h1a : _GEN_4930; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4932 = 8'h44 == _t_T_34[23:16] ? 8'h1b : _GEN_4931; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4933 = 8'h45 == _t_T_34[23:16] ? 8'h6e : _GEN_4932; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4934 = 8'h46 == _t_T_34[23:16] ? 8'h5a : _GEN_4933; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4935 = 8'h47 == _t_T_34[23:16] ? 8'ha0 : _GEN_4934; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4936 = 8'h48 == _t_T_34[23:16] ? 8'h52 : _GEN_4935; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4937 = 8'h49 == _t_T_34[23:16] ? 8'h3b : _GEN_4936; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4938 = 8'h4a == _t_T_34[23:16] ? 8'hd6 : _GEN_4937; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4939 = 8'h4b == _t_T_34[23:16] ? 8'hb3 : _GEN_4938; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4940 = 8'h4c == _t_T_34[23:16] ? 8'h29 : _GEN_4939; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4941 = 8'h4d == _t_T_34[23:16] ? 8'he3 : _GEN_4940; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4942 = 8'h4e == _t_T_34[23:16] ? 8'h2f : _GEN_4941; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4943 = 8'h4f == _t_T_34[23:16] ? 8'h84 : _GEN_4942; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4944 = 8'h50 == _t_T_34[23:16] ? 8'h53 : _GEN_4943; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4945 = 8'h51 == _t_T_34[23:16] ? 8'hd1 : _GEN_4944; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4946 = 8'h52 == _t_T_34[23:16] ? 8'h0 : _GEN_4945; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4947 = 8'h53 == _t_T_34[23:16] ? 8'hed : _GEN_4946; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4948 = 8'h54 == _t_T_34[23:16] ? 8'h20 : _GEN_4947; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4949 = 8'h55 == _t_T_34[23:16] ? 8'hfc : _GEN_4948; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4950 = 8'h56 == _t_T_34[23:16] ? 8'hb1 : _GEN_4949; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4951 = 8'h57 == _t_T_34[23:16] ? 8'h5b : _GEN_4950; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4952 = 8'h58 == _t_T_34[23:16] ? 8'h6a : _GEN_4951; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4953 = 8'h59 == _t_T_34[23:16] ? 8'hcb : _GEN_4952; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4954 = 8'h5a == _t_T_34[23:16] ? 8'hbe : _GEN_4953; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4955 = 8'h5b == _t_T_34[23:16] ? 8'h39 : _GEN_4954; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4956 = 8'h5c == _t_T_34[23:16] ? 8'h4a : _GEN_4955; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4957 = 8'h5d == _t_T_34[23:16] ? 8'h4c : _GEN_4956; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4958 = 8'h5e == _t_T_34[23:16] ? 8'h58 : _GEN_4957; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4959 = 8'h5f == _t_T_34[23:16] ? 8'hcf : _GEN_4958; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4960 = 8'h60 == _t_T_34[23:16] ? 8'hd0 : _GEN_4959; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4961 = 8'h61 == _t_T_34[23:16] ? 8'hef : _GEN_4960; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4962 = 8'h62 == _t_T_34[23:16] ? 8'haa : _GEN_4961; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4963 = 8'h63 == _t_T_34[23:16] ? 8'hfb : _GEN_4962; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4964 = 8'h64 == _t_T_34[23:16] ? 8'h43 : _GEN_4963; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4965 = 8'h65 == _t_T_34[23:16] ? 8'h4d : _GEN_4964; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4966 = 8'h66 == _t_T_34[23:16] ? 8'h33 : _GEN_4965; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4967 = 8'h67 == _t_T_34[23:16] ? 8'h85 : _GEN_4966; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4968 = 8'h68 == _t_T_34[23:16] ? 8'h45 : _GEN_4967; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4969 = 8'h69 == _t_T_34[23:16] ? 8'hf9 : _GEN_4968; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4970 = 8'h6a == _t_T_34[23:16] ? 8'h2 : _GEN_4969; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4971 = 8'h6b == _t_T_34[23:16] ? 8'h7f : _GEN_4970; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4972 = 8'h6c == _t_T_34[23:16] ? 8'h50 : _GEN_4971; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4973 = 8'h6d == _t_T_34[23:16] ? 8'h3c : _GEN_4972; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4974 = 8'h6e == _t_T_34[23:16] ? 8'h9f : _GEN_4973; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4975 = 8'h6f == _t_T_34[23:16] ? 8'ha8 : _GEN_4974; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4976 = 8'h70 == _t_T_34[23:16] ? 8'h51 : _GEN_4975; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4977 = 8'h71 == _t_T_34[23:16] ? 8'ha3 : _GEN_4976; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4978 = 8'h72 == _t_T_34[23:16] ? 8'h40 : _GEN_4977; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4979 = 8'h73 == _t_T_34[23:16] ? 8'h8f : _GEN_4978; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4980 = 8'h74 == _t_T_34[23:16] ? 8'h92 : _GEN_4979; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4981 = 8'h75 == _t_T_34[23:16] ? 8'h9d : _GEN_4980; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4982 = 8'h76 == _t_T_34[23:16] ? 8'h38 : _GEN_4981; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4983 = 8'h77 == _t_T_34[23:16] ? 8'hf5 : _GEN_4982; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4984 = 8'h78 == _t_T_34[23:16] ? 8'hbc : _GEN_4983; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4985 = 8'h79 == _t_T_34[23:16] ? 8'hb6 : _GEN_4984; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4986 = 8'h7a == _t_T_34[23:16] ? 8'hda : _GEN_4985; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4987 = 8'h7b == _t_T_34[23:16] ? 8'h21 : _GEN_4986; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4988 = 8'h7c == _t_T_34[23:16] ? 8'h10 : _GEN_4987; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4989 = 8'h7d == _t_T_34[23:16] ? 8'hff : _GEN_4988; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4990 = 8'h7e == _t_T_34[23:16] ? 8'hf3 : _GEN_4989; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4991 = 8'h7f == _t_T_34[23:16] ? 8'hd2 : _GEN_4990; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4992 = 8'h80 == _t_T_34[23:16] ? 8'hcd : _GEN_4991; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4993 = 8'h81 == _t_T_34[23:16] ? 8'hc : _GEN_4992; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4994 = 8'h82 == _t_T_34[23:16] ? 8'h13 : _GEN_4993; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4995 = 8'h83 == _t_T_34[23:16] ? 8'hec : _GEN_4994; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4996 = 8'h84 == _t_T_34[23:16] ? 8'h5f : _GEN_4995; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4997 = 8'h85 == _t_T_34[23:16] ? 8'h97 : _GEN_4996; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4998 = 8'h86 == _t_T_34[23:16] ? 8'h44 : _GEN_4997; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_4999 = 8'h87 == _t_T_34[23:16] ? 8'h17 : _GEN_4998; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5000 = 8'h88 == _t_T_34[23:16] ? 8'hc4 : _GEN_4999; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5001 = 8'h89 == _t_T_34[23:16] ? 8'ha7 : _GEN_5000; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5002 = 8'h8a == _t_T_34[23:16] ? 8'h7e : _GEN_5001; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5003 = 8'h8b == _t_T_34[23:16] ? 8'h3d : _GEN_5002; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5004 = 8'h8c == _t_T_34[23:16] ? 8'h64 : _GEN_5003; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5005 = 8'h8d == _t_T_34[23:16] ? 8'h5d : _GEN_5004; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5006 = 8'h8e == _t_T_34[23:16] ? 8'h19 : _GEN_5005; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5007 = 8'h8f == _t_T_34[23:16] ? 8'h73 : _GEN_5006; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5008 = 8'h90 == _t_T_34[23:16] ? 8'h60 : _GEN_5007; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5009 = 8'h91 == _t_T_34[23:16] ? 8'h81 : _GEN_5008; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5010 = 8'h92 == _t_T_34[23:16] ? 8'h4f : _GEN_5009; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5011 = 8'h93 == _t_T_34[23:16] ? 8'hdc : _GEN_5010; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5012 = 8'h94 == _t_T_34[23:16] ? 8'h22 : _GEN_5011; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5013 = 8'h95 == _t_T_34[23:16] ? 8'h2a : _GEN_5012; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5014 = 8'h96 == _t_T_34[23:16] ? 8'h90 : _GEN_5013; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5015 = 8'h97 == _t_T_34[23:16] ? 8'h88 : _GEN_5014; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5016 = 8'h98 == _t_T_34[23:16] ? 8'h46 : _GEN_5015; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5017 = 8'h99 == _t_T_34[23:16] ? 8'hee : _GEN_5016; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5018 = 8'h9a == _t_T_34[23:16] ? 8'hb8 : _GEN_5017; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5019 = 8'h9b == _t_T_34[23:16] ? 8'h14 : _GEN_5018; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5020 = 8'h9c == _t_T_34[23:16] ? 8'hde : _GEN_5019; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5021 = 8'h9d == _t_T_34[23:16] ? 8'h5e : _GEN_5020; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5022 = 8'h9e == _t_T_34[23:16] ? 8'hb : _GEN_5021; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5023 = 8'h9f == _t_T_34[23:16] ? 8'hdb : _GEN_5022; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5024 = 8'ha0 == _t_T_34[23:16] ? 8'he0 : _GEN_5023; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5025 = 8'ha1 == _t_T_34[23:16] ? 8'h32 : _GEN_5024; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5026 = 8'ha2 == _t_T_34[23:16] ? 8'h3a : _GEN_5025; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5027 = 8'ha3 == _t_T_34[23:16] ? 8'ha : _GEN_5026; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5028 = 8'ha4 == _t_T_34[23:16] ? 8'h49 : _GEN_5027; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5029 = 8'ha5 == _t_T_34[23:16] ? 8'h6 : _GEN_5028; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5030 = 8'ha6 == _t_T_34[23:16] ? 8'h24 : _GEN_5029; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5031 = 8'ha7 == _t_T_34[23:16] ? 8'h5c : _GEN_5030; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5032 = 8'ha8 == _t_T_34[23:16] ? 8'hc2 : _GEN_5031; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5033 = 8'ha9 == _t_T_34[23:16] ? 8'hd3 : _GEN_5032; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5034 = 8'haa == _t_T_34[23:16] ? 8'hac : _GEN_5033; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5035 = 8'hab == _t_T_34[23:16] ? 8'h62 : _GEN_5034; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5036 = 8'hac == _t_T_34[23:16] ? 8'h91 : _GEN_5035; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5037 = 8'had == _t_T_34[23:16] ? 8'h95 : _GEN_5036; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5038 = 8'hae == _t_T_34[23:16] ? 8'he4 : _GEN_5037; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5039 = 8'haf == _t_T_34[23:16] ? 8'h79 : _GEN_5038; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5040 = 8'hb0 == _t_T_34[23:16] ? 8'he7 : _GEN_5039; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5041 = 8'hb1 == _t_T_34[23:16] ? 8'hc8 : _GEN_5040; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5042 = 8'hb2 == _t_T_34[23:16] ? 8'h37 : _GEN_5041; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5043 = 8'hb3 == _t_T_34[23:16] ? 8'h6d : _GEN_5042; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5044 = 8'hb4 == _t_T_34[23:16] ? 8'h8d : _GEN_5043; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5045 = 8'hb5 == _t_T_34[23:16] ? 8'hd5 : _GEN_5044; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5046 = 8'hb6 == _t_T_34[23:16] ? 8'h4e : _GEN_5045; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5047 = 8'hb7 == _t_T_34[23:16] ? 8'ha9 : _GEN_5046; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5048 = 8'hb8 == _t_T_34[23:16] ? 8'h6c : _GEN_5047; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5049 = 8'hb9 == _t_T_34[23:16] ? 8'h56 : _GEN_5048; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5050 = 8'hba == _t_T_34[23:16] ? 8'hf4 : _GEN_5049; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5051 = 8'hbb == _t_T_34[23:16] ? 8'hea : _GEN_5050; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5052 = 8'hbc == _t_T_34[23:16] ? 8'h65 : _GEN_5051; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5053 = 8'hbd == _t_T_34[23:16] ? 8'h7a : _GEN_5052; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5054 = 8'hbe == _t_T_34[23:16] ? 8'hae : _GEN_5053; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5055 = 8'hbf == _t_T_34[23:16] ? 8'h8 : _GEN_5054; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5056 = 8'hc0 == _t_T_34[23:16] ? 8'hba : _GEN_5055; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5057 = 8'hc1 == _t_T_34[23:16] ? 8'h78 : _GEN_5056; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5058 = 8'hc2 == _t_T_34[23:16] ? 8'h25 : _GEN_5057; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5059 = 8'hc3 == _t_T_34[23:16] ? 8'h2e : _GEN_5058; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5060 = 8'hc4 == _t_T_34[23:16] ? 8'h1c : _GEN_5059; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5061 = 8'hc5 == _t_T_34[23:16] ? 8'ha6 : _GEN_5060; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5062 = 8'hc6 == _t_T_34[23:16] ? 8'hb4 : _GEN_5061; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5063 = 8'hc7 == _t_T_34[23:16] ? 8'hc6 : _GEN_5062; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5064 = 8'hc8 == _t_T_34[23:16] ? 8'he8 : _GEN_5063; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5065 = 8'hc9 == _t_T_34[23:16] ? 8'hdd : _GEN_5064; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5066 = 8'hca == _t_T_34[23:16] ? 8'h74 : _GEN_5065; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5067 = 8'hcb == _t_T_34[23:16] ? 8'h1f : _GEN_5066; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5068 = 8'hcc == _t_T_34[23:16] ? 8'h4b : _GEN_5067; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5069 = 8'hcd == _t_T_34[23:16] ? 8'hbd : _GEN_5068; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5070 = 8'hce == _t_T_34[23:16] ? 8'h8b : _GEN_5069; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5071 = 8'hcf == _t_T_34[23:16] ? 8'h8a : _GEN_5070; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5072 = 8'hd0 == _t_T_34[23:16] ? 8'h70 : _GEN_5071; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5073 = 8'hd1 == _t_T_34[23:16] ? 8'h3e : _GEN_5072; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5074 = 8'hd2 == _t_T_34[23:16] ? 8'hb5 : _GEN_5073; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5075 = 8'hd3 == _t_T_34[23:16] ? 8'h66 : _GEN_5074; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5076 = 8'hd4 == _t_T_34[23:16] ? 8'h48 : _GEN_5075; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5077 = 8'hd5 == _t_T_34[23:16] ? 8'h3 : _GEN_5076; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5078 = 8'hd6 == _t_T_34[23:16] ? 8'hf6 : _GEN_5077; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5079 = 8'hd7 == _t_T_34[23:16] ? 8'he : _GEN_5078; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5080 = 8'hd8 == _t_T_34[23:16] ? 8'h61 : _GEN_5079; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5081 = 8'hd9 == _t_T_34[23:16] ? 8'h35 : _GEN_5080; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5082 = 8'hda == _t_T_34[23:16] ? 8'h57 : _GEN_5081; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5083 = 8'hdb == _t_T_34[23:16] ? 8'hb9 : _GEN_5082; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5084 = 8'hdc == _t_T_34[23:16] ? 8'h86 : _GEN_5083; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5085 = 8'hdd == _t_T_34[23:16] ? 8'hc1 : _GEN_5084; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5086 = 8'hde == _t_T_34[23:16] ? 8'h1d : _GEN_5085; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5087 = 8'hdf == _t_T_34[23:16] ? 8'h9e : _GEN_5086; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5088 = 8'he0 == _t_T_34[23:16] ? 8'he1 : _GEN_5087; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5089 = 8'he1 == _t_T_34[23:16] ? 8'hf8 : _GEN_5088; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5090 = 8'he2 == _t_T_34[23:16] ? 8'h98 : _GEN_5089; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5091 = 8'he3 == _t_T_34[23:16] ? 8'h11 : _GEN_5090; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5092 = 8'he4 == _t_T_34[23:16] ? 8'h69 : _GEN_5091; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5093 = 8'he5 == _t_T_34[23:16] ? 8'hd9 : _GEN_5092; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5094 = 8'he6 == _t_T_34[23:16] ? 8'h8e : _GEN_5093; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5095 = 8'he7 == _t_T_34[23:16] ? 8'h94 : _GEN_5094; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5096 = 8'he8 == _t_T_34[23:16] ? 8'h9b : _GEN_5095; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5097 = 8'he9 == _t_T_34[23:16] ? 8'h1e : _GEN_5096; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5098 = 8'hea == _t_T_34[23:16] ? 8'h87 : _GEN_5097; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5099 = 8'heb == _t_T_34[23:16] ? 8'he9 : _GEN_5098; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5100 = 8'hec == _t_T_34[23:16] ? 8'hce : _GEN_5099; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5101 = 8'hed == _t_T_34[23:16] ? 8'h55 : _GEN_5100; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5102 = 8'hee == _t_T_34[23:16] ? 8'h28 : _GEN_5101; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5103 = 8'hef == _t_T_34[23:16] ? 8'hdf : _GEN_5102; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5104 = 8'hf0 == _t_T_34[23:16] ? 8'h8c : _GEN_5103; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5105 = 8'hf1 == _t_T_34[23:16] ? 8'ha1 : _GEN_5104; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5106 = 8'hf2 == _t_T_34[23:16] ? 8'h89 : _GEN_5105; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5107 = 8'hf3 == _t_T_34[23:16] ? 8'hd : _GEN_5106; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5108 = 8'hf4 == _t_T_34[23:16] ? 8'hbf : _GEN_5107; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5109 = 8'hf5 == _t_T_34[23:16] ? 8'he6 : _GEN_5108; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5110 = 8'hf6 == _t_T_34[23:16] ? 8'h42 : _GEN_5109; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5111 = 8'hf7 == _t_T_34[23:16] ? 8'h68 : _GEN_5110; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5112 = 8'hf8 == _t_T_34[23:16] ? 8'h41 : _GEN_5111; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5113 = 8'hf9 == _t_T_34[23:16] ? 8'h99 : _GEN_5112; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5114 = 8'hfa == _t_T_34[23:16] ? 8'h2d : _GEN_5113; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5115 = 8'hfb == _t_T_34[23:16] ? 8'hf : _GEN_5114; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5116 = 8'hfc == _t_T_34[23:16] ? 8'hb0 : _GEN_5115; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5117 = 8'hfd == _t_T_34[23:16] ? 8'h54 : _GEN_5116; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5118 = 8'hfe == _t_T_34[23:16] ? 8'hbb : _GEN_5117; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5119 = 8'hff == _t_T_34[23:16] ? 8'h16 : _GEN_5118; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [31:0] _t_T_39 = {_GEN_4863,_GEN_5119,_GEN_4351,_GEN_4607}; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:8]
  wire [31:0] t_4 = _t_T_39 ^ 32'h10000000; // @[src/main/scala/crypto/aes/KeySchedule.scala 59:32]
  wire [31:0] w_20 = w_16 ^ t_4; // @[src/main/scala/crypto/aes/KeySchedule.scala 63:21]
  wire [31:0] w_21 = w_17 ^ w_20; // @[src/main/scala/crypto/aes/KeySchedule.scala 63:21]
  wire [31:0] w_22 = w_18 ^ w_21; // @[src/main/scala/crypto/aes/KeySchedule.scala 63:21]
  wire [31:0] w_23 = w_19 ^ w_22; // @[src/main/scala/crypto/aes/KeySchedule.scala 63:21]
  wire [31:0] _t_T_42 = {w_23[23:0],w_23[31:24]}; // @[src/main/scala/crypto/aes/KeySchedule.scala 23:43]
  wire [7:0] _GEN_5121 = 8'h1 == _t_T_42[15:8] ? 8'h7c : 8'h63; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5122 = 8'h2 == _t_T_42[15:8] ? 8'h77 : _GEN_5121; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5123 = 8'h3 == _t_T_42[15:8] ? 8'h7b : _GEN_5122; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5124 = 8'h4 == _t_T_42[15:8] ? 8'hf2 : _GEN_5123; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5125 = 8'h5 == _t_T_42[15:8] ? 8'h6b : _GEN_5124; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5126 = 8'h6 == _t_T_42[15:8] ? 8'h6f : _GEN_5125; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5127 = 8'h7 == _t_T_42[15:8] ? 8'hc5 : _GEN_5126; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5128 = 8'h8 == _t_T_42[15:8] ? 8'h30 : _GEN_5127; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5129 = 8'h9 == _t_T_42[15:8] ? 8'h1 : _GEN_5128; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5130 = 8'ha == _t_T_42[15:8] ? 8'h67 : _GEN_5129; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5131 = 8'hb == _t_T_42[15:8] ? 8'h2b : _GEN_5130; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5132 = 8'hc == _t_T_42[15:8] ? 8'hfe : _GEN_5131; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5133 = 8'hd == _t_T_42[15:8] ? 8'hd7 : _GEN_5132; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5134 = 8'he == _t_T_42[15:8] ? 8'hab : _GEN_5133; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5135 = 8'hf == _t_T_42[15:8] ? 8'h76 : _GEN_5134; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5136 = 8'h10 == _t_T_42[15:8] ? 8'hca : _GEN_5135; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5137 = 8'h11 == _t_T_42[15:8] ? 8'h82 : _GEN_5136; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5138 = 8'h12 == _t_T_42[15:8] ? 8'hc9 : _GEN_5137; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5139 = 8'h13 == _t_T_42[15:8] ? 8'h7d : _GEN_5138; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5140 = 8'h14 == _t_T_42[15:8] ? 8'hfa : _GEN_5139; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5141 = 8'h15 == _t_T_42[15:8] ? 8'h59 : _GEN_5140; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5142 = 8'h16 == _t_T_42[15:8] ? 8'h47 : _GEN_5141; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5143 = 8'h17 == _t_T_42[15:8] ? 8'hf0 : _GEN_5142; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5144 = 8'h18 == _t_T_42[15:8] ? 8'had : _GEN_5143; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5145 = 8'h19 == _t_T_42[15:8] ? 8'hd4 : _GEN_5144; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5146 = 8'h1a == _t_T_42[15:8] ? 8'ha2 : _GEN_5145; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5147 = 8'h1b == _t_T_42[15:8] ? 8'haf : _GEN_5146; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5148 = 8'h1c == _t_T_42[15:8] ? 8'h9c : _GEN_5147; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5149 = 8'h1d == _t_T_42[15:8] ? 8'ha4 : _GEN_5148; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5150 = 8'h1e == _t_T_42[15:8] ? 8'h72 : _GEN_5149; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5151 = 8'h1f == _t_T_42[15:8] ? 8'hc0 : _GEN_5150; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5152 = 8'h20 == _t_T_42[15:8] ? 8'hb7 : _GEN_5151; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5153 = 8'h21 == _t_T_42[15:8] ? 8'hfd : _GEN_5152; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5154 = 8'h22 == _t_T_42[15:8] ? 8'h93 : _GEN_5153; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5155 = 8'h23 == _t_T_42[15:8] ? 8'h26 : _GEN_5154; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5156 = 8'h24 == _t_T_42[15:8] ? 8'h36 : _GEN_5155; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5157 = 8'h25 == _t_T_42[15:8] ? 8'h3f : _GEN_5156; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5158 = 8'h26 == _t_T_42[15:8] ? 8'hf7 : _GEN_5157; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5159 = 8'h27 == _t_T_42[15:8] ? 8'hcc : _GEN_5158; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5160 = 8'h28 == _t_T_42[15:8] ? 8'h34 : _GEN_5159; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5161 = 8'h29 == _t_T_42[15:8] ? 8'ha5 : _GEN_5160; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5162 = 8'h2a == _t_T_42[15:8] ? 8'he5 : _GEN_5161; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5163 = 8'h2b == _t_T_42[15:8] ? 8'hf1 : _GEN_5162; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5164 = 8'h2c == _t_T_42[15:8] ? 8'h71 : _GEN_5163; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5165 = 8'h2d == _t_T_42[15:8] ? 8'hd8 : _GEN_5164; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5166 = 8'h2e == _t_T_42[15:8] ? 8'h31 : _GEN_5165; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5167 = 8'h2f == _t_T_42[15:8] ? 8'h15 : _GEN_5166; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5168 = 8'h30 == _t_T_42[15:8] ? 8'h4 : _GEN_5167; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5169 = 8'h31 == _t_T_42[15:8] ? 8'hc7 : _GEN_5168; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5170 = 8'h32 == _t_T_42[15:8] ? 8'h23 : _GEN_5169; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5171 = 8'h33 == _t_T_42[15:8] ? 8'hc3 : _GEN_5170; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5172 = 8'h34 == _t_T_42[15:8] ? 8'h18 : _GEN_5171; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5173 = 8'h35 == _t_T_42[15:8] ? 8'h96 : _GEN_5172; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5174 = 8'h36 == _t_T_42[15:8] ? 8'h5 : _GEN_5173; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5175 = 8'h37 == _t_T_42[15:8] ? 8'h9a : _GEN_5174; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5176 = 8'h38 == _t_T_42[15:8] ? 8'h7 : _GEN_5175; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5177 = 8'h39 == _t_T_42[15:8] ? 8'h12 : _GEN_5176; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5178 = 8'h3a == _t_T_42[15:8] ? 8'h80 : _GEN_5177; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5179 = 8'h3b == _t_T_42[15:8] ? 8'he2 : _GEN_5178; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5180 = 8'h3c == _t_T_42[15:8] ? 8'heb : _GEN_5179; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5181 = 8'h3d == _t_T_42[15:8] ? 8'h27 : _GEN_5180; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5182 = 8'h3e == _t_T_42[15:8] ? 8'hb2 : _GEN_5181; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5183 = 8'h3f == _t_T_42[15:8] ? 8'h75 : _GEN_5182; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5184 = 8'h40 == _t_T_42[15:8] ? 8'h9 : _GEN_5183; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5185 = 8'h41 == _t_T_42[15:8] ? 8'h83 : _GEN_5184; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5186 = 8'h42 == _t_T_42[15:8] ? 8'h2c : _GEN_5185; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5187 = 8'h43 == _t_T_42[15:8] ? 8'h1a : _GEN_5186; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5188 = 8'h44 == _t_T_42[15:8] ? 8'h1b : _GEN_5187; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5189 = 8'h45 == _t_T_42[15:8] ? 8'h6e : _GEN_5188; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5190 = 8'h46 == _t_T_42[15:8] ? 8'h5a : _GEN_5189; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5191 = 8'h47 == _t_T_42[15:8] ? 8'ha0 : _GEN_5190; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5192 = 8'h48 == _t_T_42[15:8] ? 8'h52 : _GEN_5191; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5193 = 8'h49 == _t_T_42[15:8] ? 8'h3b : _GEN_5192; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5194 = 8'h4a == _t_T_42[15:8] ? 8'hd6 : _GEN_5193; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5195 = 8'h4b == _t_T_42[15:8] ? 8'hb3 : _GEN_5194; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5196 = 8'h4c == _t_T_42[15:8] ? 8'h29 : _GEN_5195; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5197 = 8'h4d == _t_T_42[15:8] ? 8'he3 : _GEN_5196; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5198 = 8'h4e == _t_T_42[15:8] ? 8'h2f : _GEN_5197; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5199 = 8'h4f == _t_T_42[15:8] ? 8'h84 : _GEN_5198; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5200 = 8'h50 == _t_T_42[15:8] ? 8'h53 : _GEN_5199; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5201 = 8'h51 == _t_T_42[15:8] ? 8'hd1 : _GEN_5200; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5202 = 8'h52 == _t_T_42[15:8] ? 8'h0 : _GEN_5201; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5203 = 8'h53 == _t_T_42[15:8] ? 8'hed : _GEN_5202; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5204 = 8'h54 == _t_T_42[15:8] ? 8'h20 : _GEN_5203; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5205 = 8'h55 == _t_T_42[15:8] ? 8'hfc : _GEN_5204; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5206 = 8'h56 == _t_T_42[15:8] ? 8'hb1 : _GEN_5205; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5207 = 8'h57 == _t_T_42[15:8] ? 8'h5b : _GEN_5206; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5208 = 8'h58 == _t_T_42[15:8] ? 8'h6a : _GEN_5207; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5209 = 8'h59 == _t_T_42[15:8] ? 8'hcb : _GEN_5208; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5210 = 8'h5a == _t_T_42[15:8] ? 8'hbe : _GEN_5209; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5211 = 8'h5b == _t_T_42[15:8] ? 8'h39 : _GEN_5210; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5212 = 8'h5c == _t_T_42[15:8] ? 8'h4a : _GEN_5211; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5213 = 8'h5d == _t_T_42[15:8] ? 8'h4c : _GEN_5212; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5214 = 8'h5e == _t_T_42[15:8] ? 8'h58 : _GEN_5213; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5215 = 8'h5f == _t_T_42[15:8] ? 8'hcf : _GEN_5214; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5216 = 8'h60 == _t_T_42[15:8] ? 8'hd0 : _GEN_5215; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5217 = 8'h61 == _t_T_42[15:8] ? 8'hef : _GEN_5216; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5218 = 8'h62 == _t_T_42[15:8] ? 8'haa : _GEN_5217; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5219 = 8'h63 == _t_T_42[15:8] ? 8'hfb : _GEN_5218; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5220 = 8'h64 == _t_T_42[15:8] ? 8'h43 : _GEN_5219; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5221 = 8'h65 == _t_T_42[15:8] ? 8'h4d : _GEN_5220; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5222 = 8'h66 == _t_T_42[15:8] ? 8'h33 : _GEN_5221; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5223 = 8'h67 == _t_T_42[15:8] ? 8'h85 : _GEN_5222; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5224 = 8'h68 == _t_T_42[15:8] ? 8'h45 : _GEN_5223; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5225 = 8'h69 == _t_T_42[15:8] ? 8'hf9 : _GEN_5224; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5226 = 8'h6a == _t_T_42[15:8] ? 8'h2 : _GEN_5225; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5227 = 8'h6b == _t_T_42[15:8] ? 8'h7f : _GEN_5226; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5228 = 8'h6c == _t_T_42[15:8] ? 8'h50 : _GEN_5227; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5229 = 8'h6d == _t_T_42[15:8] ? 8'h3c : _GEN_5228; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5230 = 8'h6e == _t_T_42[15:8] ? 8'h9f : _GEN_5229; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5231 = 8'h6f == _t_T_42[15:8] ? 8'ha8 : _GEN_5230; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5232 = 8'h70 == _t_T_42[15:8] ? 8'h51 : _GEN_5231; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5233 = 8'h71 == _t_T_42[15:8] ? 8'ha3 : _GEN_5232; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5234 = 8'h72 == _t_T_42[15:8] ? 8'h40 : _GEN_5233; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5235 = 8'h73 == _t_T_42[15:8] ? 8'h8f : _GEN_5234; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5236 = 8'h74 == _t_T_42[15:8] ? 8'h92 : _GEN_5235; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5237 = 8'h75 == _t_T_42[15:8] ? 8'h9d : _GEN_5236; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5238 = 8'h76 == _t_T_42[15:8] ? 8'h38 : _GEN_5237; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5239 = 8'h77 == _t_T_42[15:8] ? 8'hf5 : _GEN_5238; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5240 = 8'h78 == _t_T_42[15:8] ? 8'hbc : _GEN_5239; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5241 = 8'h79 == _t_T_42[15:8] ? 8'hb6 : _GEN_5240; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5242 = 8'h7a == _t_T_42[15:8] ? 8'hda : _GEN_5241; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5243 = 8'h7b == _t_T_42[15:8] ? 8'h21 : _GEN_5242; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5244 = 8'h7c == _t_T_42[15:8] ? 8'h10 : _GEN_5243; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5245 = 8'h7d == _t_T_42[15:8] ? 8'hff : _GEN_5244; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5246 = 8'h7e == _t_T_42[15:8] ? 8'hf3 : _GEN_5245; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5247 = 8'h7f == _t_T_42[15:8] ? 8'hd2 : _GEN_5246; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5248 = 8'h80 == _t_T_42[15:8] ? 8'hcd : _GEN_5247; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5249 = 8'h81 == _t_T_42[15:8] ? 8'hc : _GEN_5248; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5250 = 8'h82 == _t_T_42[15:8] ? 8'h13 : _GEN_5249; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5251 = 8'h83 == _t_T_42[15:8] ? 8'hec : _GEN_5250; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5252 = 8'h84 == _t_T_42[15:8] ? 8'h5f : _GEN_5251; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5253 = 8'h85 == _t_T_42[15:8] ? 8'h97 : _GEN_5252; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5254 = 8'h86 == _t_T_42[15:8] ? 8'h44 : _GEN_5253; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5255 = 8'h87 == _t_T_42[15:8] ? 8'h17 : _GEN_5254; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5256 = 8'h88 == _t_T_42[15:8] ? 8'hc4 : _GEN_5255; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5257 = 8'h89 == _t_T_42[15:8] ? 8'ha7 : _GEN_5256; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5258 = 8'h8a == _t_T_42[15:8] ? 8'h7e : _GEN_5257; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5259 = 8'h8b == _t_T_42[15:8] ? 8'h3d : _GEN_5258; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5260 = 8'h8c == _t_T_42[15:8] ? 8'h64 : _GEN_5259; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5261 = 8'h8d == _t_T_42[15:8] ? 8'h5d : _GEN_5260; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5262 = 8'h8e == _t_T_42[15:8] ? 8'h19 : _GEN_5261; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5263 = 8'h8f == _t_T_42[15:8] ? 8'h73 : _GEN_5262; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5264 = 8'h90 == _t_T_42[15:8] ? 8'h60 : _GEN_5263; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5265 = 8'h91 == _t_T_42[15:8] ? 8'h81 : _GEN_5264; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5266 = 8'h92 == _t_T_42[15:8] ? 8'h4f : _GEN_5265; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5267 = 8'h93 == _t_T_42[15:8] ? 8'hdc : _GEN_5266; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5268 = 8'h94 == _t_T_42[15:8] ? 8'h22 : _GEN_5267; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5269 = 8'h95 == _t_T_42[15:8] ? 8'h2a : _GEN_5268; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5270 = 8'h96 == _t_T_42[15:8] ? 8'h90 : _GEN_5269; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5271 = 8'h97 == _t_T_42[15:8] ? 8'h88 : _GEN_5270; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5272 = 8'h98 == _t_T_42[15:8] ? 8'h46 : _GEN_5271; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5273 = 8'h99 == _t_T_42[15:8] ? 8'hee : _GEN_5272; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5274 = 8'h9a == _t_T_42[15:8] ? 8'hb8 : _GEN_5273; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5275 = 8'h9b == _t_T_42[15:8] ? 8'h14 : _GEN_5274; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5276 = 8'h9c == _t_T_42[15:8] ? 8'hde : _GEN_5275; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5277 = 8'h9d == _t_T_42[15:8] ? 8'h5e : _GEN_5276; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5278 = 8'h9e == _t_T_42[15:8] ? 8'hb : _GEN_5277; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5279 = 8'h9f == _t_T_42[15:8] ? 8'hdb : _GEN_5278; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5280 = 8'ha0 == _t_T_42[15:8] ? 8'he0 : _GEN_5279; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5281 = 8'ha1 == _t_T_42[15:8] ? 8'h32 : _GEN_5280; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5282 = 8'ha2 == _t_T_42[15:8] ? 8'h3a : _GEN_5281; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5283 = 8'ha3 == _t_T_42[15:8] ? 8'ha : _GEN_5282; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5284 = 8'ha4 == _t_T_42[15:8] ? 8'h49 : _GEN_5283; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5285 = 8'ha5 == _t_T_42[15:8] ? 8'h6 : _GEN_5284; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5286 = 8'ha6 == _t_T_42[15:8] ? 8'h24 : _GEN_5285; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5287 = 8'ha7 == _t_T_42[15:8] ? 8'h5c : _GEN_5286; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5288 = 8'ha8 == _t_T_42[15:8] ? 8'hc2 : _GEN_5287; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5289 = 8'ha9 == _t_T_42[15:8] ? 8'hd3 : _GEN_5288; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5290 = 8'haa == _t_T_42[15:8] ? 8'hac : _GEN_5289; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5291 = 8'hab == _t_T_42[15:8] ? 8'h62 : _GEN_5290; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5292 = 8'hac == _t_T_42[15:8] ? 8'h91 : _GEN_5291; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5293 = 8'had == _t_T_42[15:8] ? 8'h95 : _GEN_5292; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5294 = 8'hae == _t_T_42[15:8] ? 8'he4 : _GEN_5293; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5295 = 8'haf == _t_T_42[15:8] ? 8'h79 : _GEN_5294; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5296 = 8'hb0 == _t_T_42[15:8] ? 8'he7 : _GEN_5295; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5297 = 8'hb1 == _t_T_42[15:8] ? 8'hc8 : _GEN_5296; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5298 = 8'hb2 == _t_T_42[15:8] ? 8'h37 : _GEN_5297; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5299 = 8'hb3 == _t_T_42[15:8] ? 8'h6d : _GEN_5298; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5300 = 8'hb4 == _t_T_42[15:8] ? 8'h8d : _GEN_5299; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5301 = 8'hb5 == _t_T_42[15:8] ? 8'hd5 : _GEN_5300; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5302 = 8'hb6 == _t_T_42[15:8] ? 8'h4e : _GEN_5301; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5303 = 8'hb7 == _t_T_42[15:8] ? 8'ha9 : _GEN_5302; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5304 = 8'hb8 == _t_T_42[15:8] ? 8'h6c : _GEN_5303; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5305 = 8'hb9 == _t_T_42[15:8] ? 8'h56 : _GEN_5304; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5306 = 8'hba == _t_T_42[15:8] ? 8'hf4 : _GEN_5305; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5307 = 8'hbb == _t_T_42[15:8] ? 8'hea : _GEN_5306; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5308 = 8'hbc == _t_T_42[15:8] ? 8'h65 : _GEN_5307; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5309 = 8'hbd == _t_T_42[15:8] ? 8'h7a : _GEN_5308; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5310 = 8'hbe == _t_T_42[15:8] ? 8'hae : _GEN_5309; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5311 = 8'hbf == _t_T_42[15:8] ? 8'h8 : _GEN_5310; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5312 = 8'hc0 == _t_T_42[15:8] ? 8'hba : _GEN_5311; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5313 = 8'hc1 == _t_T_42[15:8] ? 8'h78 : _GEN_5312; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5314 = 8'hc2 == _t_T_42[15:8] ? 8'h25 : _GEN_5313; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5315 = 8'hc3 == _t_T_42[15:8] ? 8'h2e : _GEN_5314; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5316 = 8'hc4 == _t_T_42[15:8] ? 8'h1c : _GEN_5315; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5317 = 8'hc5 == _t_T_42[15:8] ? 8'ha6 : _GEN_5316; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5318 = 8'hc6 == _t_T_42[15:8] ? 8'hb4 : _GEN_5317; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5319 = 8'hc7 == _t_T_42[15:8] ? 8'hc6 : _GEN_5318; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5320 = 8'hc8 == _t_T_42[15:8] ? 8'he8 : _GEN_5319; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5321 = 8'hc9 == _t_T_42[15:8] ? 8'hdd : _GEN_5320; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5322 = 8'hca == _t_T_42[15:8] ? 8'h74 : _GEN_5321; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5323 = 8'hcb == _t_T_42[15:8] ? 8'h1f : _GEN_5322; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5324 = 8'hcc == _t_T_42[15:8] ? 8'h4b : _GEN_5323; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5325 = 8'hcd == _t_T_42[15:8] ? 8'hbd : _GEN_5324; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5326 = 8'hce == _t_T_42[15:8] ? 8'h8b : _GEN_5325; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5327 = 8'hcf == _t_T_42[15:8] ? 8'h8a : _GEN_5326; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5328 = 8'hd0 == _t_T_42[15:8] ? 8'h70 : _GEN_5327; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5329 = 8'hd1 == _t_T_42[15:8] ? 8'h3e : _GEN_5328; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5330 = 8'hd2 == _t_T_42[15:8] ? 8'hb5 : _GEN_5329; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5331 = 8'hd3 == _t_T_42[15:8] ? 8'h66 : _GEN_5330; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5332 = 8'hd4 == _t_T_42[15:8] ? 8'h48 : _GEN_5331; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5333 = 8'hd5 == _t_T_42[15:8] ? 8'h3 : _GEN_5332; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5334 = 8'hd6 == _t_T_42[15:8] ? 8'hf6 : _GEN_5333; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5335 = 8'hd7 == _t_T_42[15:8] ? 8'he : _GEN_5334; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5336 = 8'hd8 == _t_T_42[15:8] ? 8'h61 : _GEN_5335; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5337 = 8'hd9 == _t_T_42[15:8] ? 8'h35 : _GEN_5336; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5338 = 8'hda == _t_T_42[15:8] ? 8'h57 : _GEN_5337; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5339 = 8'hdb == _t_T_42[15:8] ? 8'hb9 : _GEN_5338; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5340 = 8'hdc == _t_T_42[15:8] ? 8'h86 : _GEN_5339; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5341 = 8'hdd == _t_T_42[15:8] ? 8'hc1 : _GEN_5340; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5342 = 8'hde == _t_T_42[15:8] ? 8'h1d : _GEN_5341; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5343 = 8'hdf == _t_T_42[15:8] ? 8'h9e : _GEN_5342; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5344 = 8'he0 == _t_T_42[15:8] ? 8'he1 : _GEN_5343; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5345 = 8'he1 == _t_T_42[15:8] ? 8'hf8 : _GEN_5344; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5346 = 8'he2 == _t_T_42[15:8] ? 8'h98 : _GEN_5345; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5347 = 8'he3 == _t_T_42[15:8] ? 8'h11 : _GEN_5346; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5348 = 8'he4 == _t_T_42[15:8] ? 8'h69 : _GEN_5347; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5349 = 8'he5 == _t_T_42[15:8] ? 8'hd9 : _GEN_5348; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5350 = 8'he6 == _t_T_42[15:8] ? 8'h8e : _GEN_5349; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5351 = 8'he7 == _t_T_42[15:8] ? 8'h94 : _GEN_5350; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5352 = 8'he8 == _t_T_42[15:8] ? 8'h9b : _GEN_5351; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5353 = 8'he9 == _t_T_42[15:8] ? 8'h1e : _GEN_5352; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5354 = 8'hea == _t_T_42[15:8] ? 8'h87 : _GEN_5353; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5355 = 8'heb == _t_T_42[15:8] ? 8'he9 : _GEN_5354; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5356 = 8'hec == _t_T_42[15:8] ? 8'hce : _GEN_5355; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5357 = 8'hed == _t_T_42[15:8] ? 8'h55 : _GEN_5356; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5358 = 8'hee == _t_T_42[15:8] ? 8'h28 : _GEN_5357; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5359 = 8'hef == _t_T_42[15:8] ? 8'hdf : _GEN_5358; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5360 = 8'hf0 == _t_T_42[15:8] ? 8'h8c : _GEN_5359; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5361 = 8'hf1 == _t_T_42[15:8] ? 8'ha1 : _GEN_5360; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5362 = 8'hf2 == _t_T_42[15:8] ? 8'h89 : _GEN_5361; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5363 = 8'hf3 == _t_T_42[15:8] ? 8'hd : _GEN_5362; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5364 = 8'hf4 == _t_T_42[15:8] ? 8'hbf : _GEN_5363; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5365 = 8'hf5 == _t_T_42[15:8] ? 8'he6 : _GEN_5364; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5366 = 8'hf6 == _t_T_42[15:8] ? 8'h42 : _GEN_5365; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5367 = 8'hf7 == _t_T_42[15:8] ? 8'h68 : _GEN_5366; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5368 = 8'hf8 == _t_T_42[15:8] ? 8'h41 : _GEN_5367; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5369 = 8'hf9 == _t_T_42[15:8] ? 8'h99 : _GEN_5368; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5370 = 8'hfa == _t_T_42[15:8] ? 8'h2d : _GEN_5369; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5371 = 8'hfb == _t_T_42[15:8] ? 8'hf : _GEN_5370; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5372 = 8'hfc == _t_T_42[15:8] ? 8'hb0 : _GEN_5371; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5373 = 8'hfd == _t_T_42[15:8] ? 8'h54 : _GEN_5372; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5374 = 8'hfe == _t_T_42[15:8] ? 8'hbb : _GEN_5373; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5375 = 8'hff == _t_T_42[15:8] ? 8'h16 : _GEN_5374; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5377 = 8'h1 == _t_T_42[7:0] ? 8'h7c : 8'h63; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5378 = 8'h2 == _t_T_42[7:0] ? 8'h77 : _GEN_5377; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5379 = 8'h3 == _t_T_42[7:0] ? 8'h7b : _GEN_5378; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5380 = 8'h4 == _t_T_42[7:0] ? 8'hf2 : _GEN_5379; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5381 = 8'h5 == _t_T_42[7:0] ? 8'h6b : _GEN_5380; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5382 = 8'h6 == _t_T_42[7:0] ? 8'h6f : _GEN_5381; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5383 = 8'h7 == _t_T_42[7:0] ? 8'hc5 : _GEN_5382; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5384 = 8'h8 == _t_T_42[7:0] ? 8'h30 : _GEN_5383; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5385 = 8'h9 == _t_T_42[7:0] ? 8'h1 : _GEN_5384; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5386 = 8'ha == _t_T_42[7:0] ? 8'h67 : _GEN_5385; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5387 = 8'hb == _t_T_42[7:0] ? 8'h2b : _GEN_5386; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5388 = 8'hc == _t_T_42[7:0] ? 8'hfe : _GEN_5387; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5389 = 8'hd == _t_T_42[7:0] ? 8'hd7 : _GEN_5388; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5390 = 8'he == _t_T_42[7:0] ? 8'hab : _GEN_5389; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5391 = 8'hf == _t_T_42[7:0] ? 8'h76 : _GEN_5390; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5392 = 8'h10 == _t_T_42[7:0] ? 8'hca : _GEN_5391; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5393 = 8'h11 == _t_T_42[7:0] ? 8'h82 : _GEN_5392; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5394 = 8'h12 == _t_T_42[7:0] ? 8'hc9 : _GEN_5393; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5395 = 8'h13 == _t_T_42[7:0] ? 8'h7d : _GEN_5394; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5396 = 8'h14 == _t_T_42[7:0] ? 8'hfa : _GEN_5395; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5397 = 8'h15 == _t_T_42[7:0] ? 8'h59 : _GEN_5396; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5398 = 8'h16 == _t_T_42[7:0] ? 8'h47 : _GEN_5397; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5399 = 8'h17 == _t_T_42[7:0] ? 8'hf0 : _GEN_5398; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5400 = 8'h18 == _t_T_42[7:0] ? 8'had : _GEN_5399; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5401 = 8'h19 == _t_T_42[7:0] ? 8'hd4 : _GEN_5400; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5402 = 8'h1a == _t_T_42[7:0] ? 8'ha2 : _GEN_5401; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5403 = 8'h1b == _t_T_42[7:0] ? 8'haf : _GEN_5402; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5404 = 8'h1c == _t_T_42[7:0] ? 8'h9c : _GEN_5403; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5405 = 8'h1d == _t_T_42[7:0] ? 8'ha4 : _GEN_5404; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5406 = 8'h1e == _t_T_42[7:0] ? 8'h72 : _GEN_5405; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5407 = 8'h1f == _t_T_42[7:0] ? 8'hc0 : _GEN_5406; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5408 = 8'h20 == _t_T_42[7:0] ? 8'hb7 : _GEN_5407; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5409 = 8'h21 == _t_T_42[7:0] ? 8'hfd : _GEN_5408; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5410 = 8'h22 == _t_T_42[7:0] ? 8'h93 : _GEN_5409; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5411 = 8'h23 == _t_T_42[7:0] ? 8'h26 : _GEN_5410; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5412 = 8'h24 == _t_T_42[7:0] ? 8'h36 : _GEN_5411; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5413 = 8'h25 == _t_T_42[7:0] ? 8'h3f : _GEN_5412; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5414 = 8'h26 == _t_T_42[7:0] ? 8'hf7 : _GEN_5413; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5415 = 8'h27 == _t_T_42[7:0] ? 8'hcc : _GEN_5414; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5416 = 8'h28 == _t_T_42[7:0] ? 8'h34 : _GEN_5415; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5417 = 8'h29 == _t_T_42[7:0] ? 8'ha5 : _GEN_5416; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5418 = 8'h2a == _t_T_42[7:0] ? 8'he5 : _GEN_5417; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5419 = 8'h2b == _t_T_42[7:0] ? 8'hf1 : _GEN_5418; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5420 = 8'h2c == _t_T_42[7:0] ? 8'h71 : _GEN_5419; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5421 = 8'h2d == _t_T_42[7:0] ? 8'hd8 : _GEN_5420; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5422 = 8'h2e == _t_T_42[7:0] ? 8'h31 : _GEN_5421; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5423 = 8'h2f == _t_T_42[7:0] ? 8'h15 : _GEN_5422; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5424 = 8'h30 == _t_T_42[7:0] ? 8'h4 : _GEN_5423; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5425 = 8'h31 == _t_T_42[7:0] ? 8'hc7 : _GEN_5424; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5426 = 8'h32 == _t_T_42[7:0] ? 8'h23 : _GEN_5425; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5427 = 8'h33 == _t_T_42[7:0] ? 8'hc3 : _GEN_5426; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5428 = 8'h34 == _t_T_42[7:0] ? 8'h18 : _GEN_5427; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5429 = 8'h35 == _t_T_42[7:0] ? 8'h96 : _GEN_5428; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5430 = 8'h36 == _t_T_42[7:0] ? 8'h5 : _GEN_5429; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5431 = 8'h37 == _t_T_42[7:0] ? 8'h9a : _GEN_5430; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5432 = 8'h38 == _t_T_42[7:0] ? 8'h7 : _GEN_5431; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5433 = 8'h39 == _t_T_42[7:0] ? 8'h12 : _GEN_5432; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5434 = 8'h3a == _t_T_42[7:0] ? 8'h80 : _GEN_5433; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5435 = 8'h3b == _t_T_42[7:0] ? 8'he2 : _GEN_5434; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5436 = 8'h3c == _t_T_42[7:0] ? 8'heb : _GEN_5435; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5437 = 8'h3d == _t_T_42[7:0] ? 8'h27 : _GEN_5436; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5438 = 8'h3e == _t_T_42[7:0] ? 8'hb2 : _GEN_5437; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5439 = 8'h3f == _t_T_42[7:0] ? 8'h75 : _GEN_5438; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5440 = 8'h40 == _t_T_42[7:0] ? 8'h9 : _GEN_5439; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5441 = 8'h41 == _t_T_42[7:0] ? 8'h83 : _GEN_5440; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5442 = 8'h42 == _t_T_42[7:0] ? 8'h2c : _GEN_5441; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5443 = 8'h43 == _t_T_42[7:0] ? 8'h1a : _GEN_5442; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5444 = 8'h44 == _t_T_42[7:0] ? 8'h1b : _GEN_5443; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5445 = 8'h45 == _t_T_42[7:0] ? 8'h6e : _GEN_5444; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5446 = 8'h46 == _t_T_42[7:0] ? 8'h5a : _GEN_5445; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5447 = 8'h47 == _t_T_42[7:0] ? 8'ha0 : _GEN_5446; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5448 = 8'h48 == _t_T_42[7:0] ? 8'h52 : _GEN_5447; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5449 = 8'h49 == _t_T_42[7:0] ? 8'h3b : _GEN_5448; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5450 = 8'h4a == _t_T_42[7:0] ? 8'hd6 : _GEN_5449; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5451 = 8'h4b == _t_T_42[7:0] ? 8'hb3 : _GEN_5450; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5452 = 8'h4c == _t_T_42[7:0] ? 8'h29 : _GEN_5451; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5453 = 8'h4d == _t_T_42[7:0] ? 8'he3 : _GEN_5452; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5454 = 8'h4e == _t_T_42[7:0] ? 8'h2f : _GEN_5453; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5455 = 8'h4f == _t_T_42[7:0] ? 8'h84 : _GEN_5454; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5456 = 8'h50 == _t_T_42[7:0] ? 8'h53 : _GEN_5455; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5457 = 8'h51 == _t_T_42[7:0] ? 8'hd1 : _GEN_5456; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5458 = 8'h52 == _t_T_42[7:0] ? 8'h0 : _GEN_5457; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5459 = 8'h53 == _t_T_42[7:0] ? 8'hed : _GEN_5458; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5460 = 8'h54 == _t_T_42[7:0] ? 8'h20 : _GEN_5459; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5461 = 8'h55 == _t_T_42[7:0] ? 8'hfc : _GEN_5460; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5462 = 8'h56 == _t_T_42[7:0] ? 8'hb1 : _GEN_5461; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5463 = 8'h57 == _t_T_42[7:0] ? 8'h5b : _GEN_5462; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5464 = 8'h58 == _t_T_42[7:0] ? 8'h6a : _GEN_5463; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5465 = 8'h59 == _t_T_42[7:0] ? 8'hcb : _GEN_5464; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5466 = 8'h5a == _t_T_42[7:0] ? 8'hbe : _GEN_5465; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5467 = 8'h5b == _t_T_42[7:0] ? 8'h39 : _GEN_5466; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5468 = 8'h5c == _t_T_42[7:0] ? 8'h4a : _GEN_5467; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5469 = 8'h5d == _t_T_42[7:0] ? 8'h4c : _GEN_5468; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5470 = 8'h5e == _t_T_42[7:0] ? 8'h58 : _GEN_5469; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5471 = 8'h5f == _t_T_42[7:0] ? 8'hcf : _GEN_5470; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5472 = 8'h60 == _t_T_42[7:0] ? 8'hd0 : _GEN_5471; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5473 = 8'h61 == _t_T_42[7:0] ? 8'hef : _GEN_5472; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5474 = 8'h62 == _t_T_42[7:0] ? 8'haa : _GEN_5473; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5475 = 8'h63 == _t_T_42[7:0] ? 8'hfb : _GEN_5474; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5476 = 8'h64 == _t_T_42[7:0] ? 8'h43 : _GEN_5475; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5477 = 8'h65 == _t_T_42[7:0] ? 8'h4d : _GEN_5476; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5478 = 8'h66 == _t_T_42[7:0] ? 8'h33 : _GEN_5477; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5479 = 8'h67 == _t_T_42[7:0] ? 8'h85 : _GEN_5478; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5480 = 8'h68 == _t_T_42[7:0] ? 8'h45 : _GEN_5479; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5481 = 8'h69 == _t_T_42[7:0] ? 8'hf9 : _GEN_5480; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5482 = 8'h6a == _t_T_42[7:0] ? 8'h2 : _GEN_5481; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5483 = 8'h6b == _t_T_42[7:0] ? 8'h7f : _GEN_5482; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5484 = 8'h6c == _t_T_42[7:0] ? 8'h50 : _GEN_5483; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5485 = 8'h6d == _t_T_42[7:0] ? 8'h3c : _GEN_5484; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5486 = 8'h6e == _t_T_42[7:0] ? 8'h9f : _GEN_5485; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5487 = 8'h6f == _t_T_42[7:0] ? 8'ha8 : _GEN_5486; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5488 = 8'h70 == _t_T_42[7:0] ? 8'h51 : _GEN_5487; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5489 = 8'h71 == _t_T_42[7:0] ? 8'ha3 : _GEN_5488; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5490 = 8'h72 == _t_T_42[7:0] ? 8'h40 : _GEN_5489; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5491 = 8'h73 == _t_T_42[7:0] ? 8'h8f : _GEN_5490; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5492 = 8'h74 == _t_T_42[7:0] ? 8'h92 : _GEN_5491; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5493 = 8'h75 == _t_T_42[7:0] ? 8'h9d : _GEN_5492; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5494 = 8'h76 == _t_T_42[7:0] ? 8'h38 : _GEN_5493; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5495 = 8'h77 == _t_T_42[7:0] ? 8'hf5 : _GEN_5494; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5496 = 8'h78 == _t_T_42[7:0] ? 8'hbc : _GEN_5495; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5497 = 8'h79 == _t_T_42[7:0] ? 8'hb6 : _GEN_5496; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5498 = 8'h7a == _t_T_42[7:0] ? 8'hda : _GEN_5497; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5499 = 8'h7b == _t_T_42[7:0] ? 8'h21 : _GEN_5498; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5500 = 8'h7c == _t_T_42[7:0] ? 8'h10 : _GEN_5499; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5501 = 8'h7d == _t_T_42[7:0] ? 8'hff : _GEN_5500; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5502 = 8'h7e == _t_T_42[7:0] ? 8'hf3 : _GEN_5501; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5503 = 8'h7f == _t_T_42[7:0] ? 8'hd2 : _GEN_5502; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5504 = 8'h80 == _t_T_42[7:0] ? 8'hcd : _GEN_5503; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5505 = 8'h81 == _t_T_42[7:0] ? 8'hc : _GEN_5504; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5506 = 8'h82 == _t_T_42[7:0] ? 8'h13 : _GEN_5505; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5507 = 8'h83 == _t_T_42[7:0] ? 8'hec : _GEN_5506; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5508 = 8'h84 == _t_T_42[7:0] ? 8'h5f : _GEN_5507; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5509 = 8'h85 == _t_T_42[7:0] ? 8'h97 : _GEN_5508; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5510 = 8'h86 == _t_T_42[7:0] ? 8'h44 : _GEN_5509; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5511 = 8'h87 == _t_T_42[7:0] ? 8'h17 : _GEN_5510; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5512 = 8'h88 == _t_T_42[7:0] ? 8'hc4 : _GEN_5511; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5513 = 8'h89 == _t_T_42[7:0] ? 8'ha7 : _GEN_5512; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5514 = 8'h8a == _t_T_42[7:0] ? 8'h7e : _GEN_5513; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5515 = 8'h8b == _t_T_42[7:0] ? 8'h3d : _GEN_5514; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5516 = 8'h8c == _t_T_42[7:0] ? 8'h64 : _GEN_5515; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5517 = 8'h8d == _t_T_42[7:0] ? 8'h5d : _GEN_5516; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5518 = 8'h8e == _t_T_42[7:0] ? 8'h19 : _GEN_5517; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5519 = 8'h8f == _t_T_42[7:0] ? 8'h73 : _GEN_5518; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5520 = 8'h90 == _t_T_42[7:0] ? 8'h60 : _GEN_5519; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5521 = 8'h91 == _t_T_42[7:0] ? 8'h81 : _GEN_5520; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5522 = 8'h92 == _t_T_42[7:0] ? 8'h4f : _GEN_5521; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5523 = 8'h93 == _t_T_42[7:0] ? 8'hdc : _GEN_5522; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5524 = 8'h94 == _t_T_42[7:0] ? 8'h22 : _GEN_5523; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5525 = 8'h95 == _t_T_42[7:0] ? 8'h2a : _GEN_5524; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5526 = 8'h96 == _t_T_42[7:0] ? 8'h90 : _GEN_5525; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5527 = 8'h97 == _t_T_42[7:0] ? 8'h88 : _GEN_5526; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5528 = 8'h98 == _t_T_42[7:0] ? 8'h46 : _GEN_5527; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5529 = 8'h99 == _t_T_42[7:0] ? 8'hee : _GEN_5528; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5530 = 8'h9a == _t_T_42[7:0] ? 8'hb8 : _GEN_5529; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5531 = 8'h9b == _t_T_42[7:0] ? 8'h14 : _GEN_5530; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5532 = 8'h9c == _t_T_42[7:0] ? 8'hde : _GEN_5531; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5533 = 8'h9d == _t_T_42[7:0] ? 8'h5e : _GEN_5532; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5534 = 8'h9e == _t_T_42[7:0] ? 8'hb : _GEN_5533; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5535 = 8'h9f == _t_T_42[7:0] ? 8'hdb : _GEN_5534; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5536 = 8'ha0 == _t_T_42[7:0] ? 8'he0 : _GEN_5535; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5537 = 8'ha1 == _t_T_42[7:0] ? 8'h32 : _GEN_5536; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5538 = 8'ha2 == _t_T_42[7:0] ? 8'h3a : _GEN_5537; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5539 = 8'ha3 == _t_T_42[7:0] ? 8'ha : _GEN_5538; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5540 = 8'ha4 == _t_T_42[7:0] ? 8'h49 : _GEN_5539; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5541 = 8'ha5 == _t_T_42[7:0] ? 8'h6 : _GEN_5540; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5542 = 8'ha6 == _t_T_42[7:0] ? 8'h24 : _GEN_5541; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5543 = 8'ha7 == _t_T_42[7:0] ? 8'h5c : _GEN_5542; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5544 = 8'ha8 == _t_T_42[7:0] ? 8'hc2 : _GEN_5543; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5545 = 8'ha9 == _t_T_42[7:0] ? 8'hd3 : _GEN_5544; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5546 = 8'haa == _t_T_42[7:0] ? 8'hac : _GEN_5545; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5547 = 8'hab == _t_T_42[7:0] ? 8'h62 : _GEN_5546; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5548 = 8'hac == _t_T_42[7:0] ? 8'h91 : _GEN_5547; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5549 = 8'had == _t_T_42[7:0] ? 8'h95 : _GEN_5548; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5550 = 8'hae == _t_T_42[7:0] ? 8'he4 : _GEN_5549; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5551 = 8'haf == _t_T_42[7:0] ? 8'h79 : _GEN_5550; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5552 = 8'hb0 == _t_T_42[7:0] ? 8'he7 : _GEN_5551; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5553 = 8'hb1 == _t_T_42[7:0] ? 8'hc8 : _GEN_5552; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5554 = 8'hb2 == _t_T_42[7:0] ? 8'h37 : _GEN_5553; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5555 = 8'hb3 == _t_T_42[7:0] ? 8'h6d : _GEN_5554; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5556 = 8'hb4 == _t_T_42[7:0] ? 8'h8d : _GEN_5555; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5557 = 8'hb5 == _t_T_42[7:0] ? 8'hd5 : _GEN_5556; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5558 = 8'hb6 == _t_T_42[7:0] ? 8'h4e : _GEN_5557; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5559 = 8'hb7 == _t_T_42[7:0] ? 8'ha9 : _GEN_5558; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5560 = 8'hb8 == _t_T_42[7:0] ? 8'h6c : _GEN_5559; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5561 = 8'hb9 == _t_T_42[7:0] ? 8'h56 : _GEN_5560; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5562 = 8'hba == _t_T_42[7:0] ? 8'hf4 : _GEN_5561; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5563 = 8'hbb == _t_T_42[7:0] ? 8'hea : _GEN_5562; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5564 = 8'hbc == _t_T_42[7:0] ? 8'h65 : _GEN_5563; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5565 = 8'hbd == _t_T_42[7:0] ? 8'h7a : _GEN_5564; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5566 = 8'hbe == _t_T_42[7:0] ? 8'hae : _GEN_5565; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5567 = 8'hbf == _t_T_42[7:0] ? 8'h8 : _GEN_5566; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5568 = 8'hc0 == _t_T_42[7:0] ? 8'hba : _GEN_5567; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5569 = 8'hc1 == _t_T_42[7:0] ? 8'h78 : _GEN_5568; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5570 = 8'hc2 == _t_T_42[7:0] ? 8'h25 : _GEN_5569; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5571 = 8'hc3 == _t_T_42[7:0] ? 8'h2e : _GEN_5570; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5572 = 8'hc4 == _t_T_42[7:0] ? 8'h1c : _GEN_5571; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5573 = 8'hc5 == _t_T_42[7:0] ? 8'ha6 : _GEN_5572; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5574 = 8'hc6 == _t_T_42[7:0] ? 8'hb4 : _GEN_5573; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5575 = 8'hc7 == _t_T_42[7:0] ? 8'hc6 : _GEN_5574; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5576 = 8'hc8 == _t_T_42[7:0] ? 8'he8 : _GEN_5575; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5577 = 8'hc9 == _t_T_42[7:0] ? 8'hdd : _GEN_5576; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5578 = 8'hca == _t_T_42[7:0] ? 8'h74 : _GEN_5577; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5579 = 8'hcb == _t_T_42[7:0] ? 8'h1f : _GEN_5578; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5580 = 8'hcc == _t_T_42[7:0] ? 8'h4b : _GEN_5579; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5581 = 8'hcd == _t_T_42[7:0] ? 8'hbd : _GEN_5580; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5582 = 8'hce == _t_T_42[7:0] ? 8'h8b : _GEN_5581; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5583 = 8'hcf == _t_T_42[7:0] ? 8'h8a : _GEN_5582; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5584 = 8'hd0 == _t_T_42[7:0] ? 8'h70 : _GEN_5583; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5585 = 8'hd1 == _t_T_42[7:0] ? 8'h3e : _GEN_5584; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5586 = 8'hd2 == _t_T_42[7:0] ? 8'hb5 : _GEN_5585; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5587 = 8'hd3 == _t_T_42[7:0] ? 8'h66 : _GEN_5586; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5588 = 8'hd4 == _t_T_42[7:0] ? 8'h48 : _GEN_5587; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5589 = 8'hd5 == _t_T_42[7:0] ? 8'h3 : _GEN_5588; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5590 = 8'hd6 == _t_T_42[7:0] ? 8'hf6 : _GEN_5589; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5591 = 8'hd7 == _t_T_42[7:0] ? 8'he : _GEN_5590; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5592 = 8'hd8 == _t_T_42[7:0] ? 8'h61 : _GEN_5591; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5593 = 8'hd9 == _t_T_42[7:0] ? 8'h35 : _GEN_5592; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5594 = 8'hda == _t_T_42[7:0] ? 8'h57 : _GEN_5593; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5595 = 8'hdb == _t_T_42[7:0] ? 8'hb9 : _GEN_5594; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5596 = 8'hdc == _t_T_42[7:0] ? 8'h86 : _GEN_5595; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5597 = 8'hdd == _t_T_42[7:0] ? 8'hc1 : _GEN_5596; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5598 = 8'hde == _t_T_42[7:0] ? 8'h1d : _GEN_5597; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5599 = 8'hdf == _t_T_42[7:0] ? 8'h9e : _GEN_5598; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5600 = 8'he0 == _t_T_42[7:0] ? 8'he1 : _GEN_5599; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5601 = 8'he1 == _t_T_42[7:0] ? 8'hf8 : _GEN_5600; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5602 = 8'he2 == _t_T_42[7:0] ? 8'h98 : _GEN_5601; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5603 = 8'he3 == _t_T_42[7:0] ? 8'h11 : _GEN_5602; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5604 = 8'he4 == _t_T_42[7:0] ? 8'h69 : _GEN_5603; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5605 = 8'he5 == _t_T_42[7:0] ? 8'hd9 : _GEN_5604; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5606 = 8'he6 == _t_T_42[7:0] ? 8'h8e : _GEN_5605; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5607 = 8'he7 == _t_T_42[7:0] ? 8'h94 : _GEN_5606; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5608 = 8'he8 == _t_T_42[7:0] ? 8'h9b : _GEN_5607; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5609 = 8'he9 == _t_T_42[7:0] ? 8'h1e : _GEN_5608; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5610 = 8'hea == _t_T_42[7:0] ? 8'h87 : _GEN_5609; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5611 = 8'heb == _t_T_42[7:0] ? 8'he9 : _GEN_5610; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5612 = 8'hec == _t_T_42[7:0] ? 8'hce : _GEN_5611; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5613 = 8'hed == _t_T_42[7:0] ? 8'h55 : _GEN_5612; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5614 = 8'hee == _t_T_42[7:0] ? 8'h28 : _GEN_5613; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5615 = 8'hef == _t_T_42[7:0] ? 8'hdf : _GEN_5614; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5616 = 8'hf0 == _t_T_42[7:0] ? 8'h8c : _GEN_5615; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5617 = 8'hf1 == _t_T_42[7:0] ? 8'ha1 : _GEN_5616; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5618 = 8'hf2 == _t_T_42[7:0] ? 8'h89 : _GEN_5617; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5619 = 8'hf3 == _t_T_42[7:0] ? 8'hd : _GEN_5618; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5620 = 8'hf4 == _t_T_42[7:0] ? 8'hbf : _GEN_5619; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5621 = 8'hf5 == _t_T_42[7:0] ? 8'he6 : _GEN_5620; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5622 = 8'hf6 == _t_T_42[7:0] ? 8'h42 : _GEN_5621; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5623 = 8'hf7 == _t_T_42[7:0] ? 8'h68 : _GEN_5622; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5624 = 8'hf8 == _t_T_42[7:0] ? 8'h41 : _GEN_5623; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5625 = 8'hf9 == _t_T_42[7:0] ? 8'h99 : _GEN_5624; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5626 = 8'hfa == _t_T_42[7:0] ? 8'h2d : _GEN_5625; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5627 = 8'hfb == _t_T_42[7:0] ? 8'hf : _GEN_5626; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5628 = 8'hfc == _t_T_42[7:0] ? 8'hb0 : _GEN_5627; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5629 = 8'hfd == _t_T_42[7:0] ? 8'h54 : _GEN_5628; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5630 = 8'hfe == _t_T_42[7:0] ? 8'hbb : _GEN_5629; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5631 = 8'hff == _t_T_42[7:0] ? 8'h16 : _GEN_5630; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5633 = 8'h1 == _t_T_42[31:24] ? 8'h7c : 8'h63; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5634 = 8'h2 == _t_T_42[31:24] ? 8'h77 : _GEN_5633; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5635 = 8'h3 == _t_T_42[31:24] ? 8'h7b : _GEN_5634; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5636 = 8'h4 == _t_T_42[31:24] ? 8'hf2 : _GEN_5635; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5637 = 8'h5 == _t_T_42[31:24] ? 8'h6b : _GEN_5636; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5638 = 8'h6 == _t_T_42[31:24] ? 8'h6f : _GEN_5637; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5639 = 8'h7 == _t_T_42[31:24] ? 8'hc5 : _GEN_5638; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5640 = 8'h8 == _t_T_42[31:24] ? 8'h30 : _GEN_5639; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5641 = 8'h9 == _t_T_42[31:24] ? 8'h1 : _GEN_5640; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5642 = 8'ha == _t_T_42[31:24] ? 8'h67 : _GEN_5641; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5643 = 8'hb == _t_T_42[31:24] ? 8'h2b : _GEN_5642; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5644 = 8'hc == _t_T_42[31:24] ? 8'hfe : _GEN_5643; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5645 = 8'hd == _t_T_42[31:24] ? 8'hd7 : _GEN_5644; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5646 = 8'he == _t_T_42[31:24] ? 8'hab : _GEN_5645; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5647 = 8'hf == _t_T_42[31:24] ? 8'h76 : _GEN_5646; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5648 = 8'h10 == _t_T_42[31:24] ? 8'hca : _GEN_5647; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5649 = 8'h11 == _t_T_42[31:24] ? 8'h82 : _GEN_5648; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5650 = 8'h12 == _t_T_42[31:24] ? 8'hc9 : _GEN_5649; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5651 = 8'h13 == _t_T_42[31:24] ? 8'h7d : _GEN_5650; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5652 = 8'h14 == _t_T_42[31:24] ? 8'hfa : _GEN_5651; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5653 = 8'h15 == _t_T_42[31:24] ? 8'h59 : _GEN_5652; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5654 = 8'h16 == _t_T_42[31:24] ? 8'h47 : _GEN_5653; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5655 = 8'h17 == _t_T_42[31:24] ? 8'hf0 : _GEN_5654; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5656 = 8'h18 == _t_T_42[31:24] ? 8'had : _GEN_5655; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5657 = 8'h19 == _t_T_42[31:24] ? 8'hd4 : _GEN_5656; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5658 = 8'h1a == _t_T_42[31:24] ? 8'ha2 : _GEN_5657; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5659 = 8'h1b == _t_T_42[31:24] ? 8'haf : _GEN_5658; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5660 = 8'h1c == _t_T_42[31:24] ? 8'h9c : _GEN_5659; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5661 = 8'h1d == _t_T_42[31:24] ? 8'ha4 : _GEN_5660; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5662 = 8'h1e == _t_T_42[31:24] ? 8'h72 : _GEN_5661; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5663 = 8'h1f == _t_T_42[31:24] ? 8'hc0 : _GEN_5662; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5664 = 8'h20 == _t_T_42[31:24] ? 8'hb7 : _GEN_5663; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5665 = 8'h21 == _t_T_42[31:24] ? 8'hfd : _GEN_5664; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5666 = 8'h22 == _t_T_42[31:24] ? 8'h93 : _GEN_5665; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5667 = 8'h23 == _t_T_42[31:24] ? 8'h26 : _GEN_5666; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5668 = 8'h24 == _t_T_42[31:24] ? 8'h36 : _GEN_5667; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5669 = 8'h25 == _t_T_42[31:24] ? 8'h3f : _GEN_5668; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5670 = 8'h26 == _t_T_42[31:24] ? 8'hf7 : _GEN_5669; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5671 = 8'h27 == _t_T_42[31:24] ? 8'hcc : _GEN_5670; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5672 = 8'h28 == _t_T_42[31:24] ? 8'h34 : _GEN_5671; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5673 = 8'h29 == _t_T_42[31:24] ? 8'ha5 : _GEN_5672; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5674 = 8'h2a == _t_T_42[31:24] ? 8'he5 : _GEN_5673; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5675 = 8'h2b == _t_T_42[31:24] ? 8'hf1 : _GEN_5674; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5676 = 8'h2c == _t_T_42[31:24] ? 8'h71 : _GEN_5675; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5677 = 8'h2d == _t_T_42[31:24] ? 8'hd8 : _GEN_5676; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5678 = 8'h2e == _t_T_42[31:24] ? 8'h31 : _GEN_5677; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5679 = 8'h2f == _t_T_42[31:24] ? 8'h15 : _GEN_5678; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5680 = 8'h30 == _t_T_42[31:24] ? 8'h4 : _GEN_5679; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5681 = 8'h31 == _t_T_42[31:24] ? 8'hc7 : _GEN_5680; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5682 = 8'h32 == _t_T_42[31:24] ? 8'h23 : _GEN_5681; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5683 = 8'h33 == _t_T_42[31:24] ? 8'hc3 : _GEN_5682; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5684 = 8'h34 == _t_T_42[31:24] ? 8'h18 : _GEN_5683; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5685 = 8'h35 == _t_T_42[31:24] ? 8'h96 : _GEN_5684; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5686 = 8'h36 == _t_T_42[31:24] ? 8'h5 : _GEN_5685; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5687 = 8'h37 == _t_T_42[31:24] ? 8'h9a : _GEN_5686; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5688 = 8'h38 == _t_T_42[31:24] ? 8'h7 : _GEN_5687; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5689 = 8'h39 == _t_T_42[31:24] ? 8'h12 : _GEN_5688; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5690 = 8'h3a == _t_T_42[31:24] ? 8'h80 : _GEN_5689; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5691 = 8'h3b == _t_T_42[31:24] ? 8'he2 : _GEN_5690; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5692 = 8'h3c == _t_T_42[31:24] ? 8'heb : _GEN_5691; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5693 = 8'h3d == _t_T_42[31:24] ? 8'h27 : _GEN_5692; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5694 = 8'h3e == _t_T_42[31:24] ? 8'hb2 : _GEN_5693; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5695 = 8'h3f == _t_T_42[31:24] ? 8'h75 : _GEN_5694; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5696 = 8'h40 == _t_T_42[31:24] ? 8'h9 : _GEN_5695; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5697 = 8'h41 == _t_T_42[31:24] ? 8'h83 : _GEN_5696; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5698 = 8'h42 == _t_T_42[31:24] ? 8'h2c : _GEN_5697; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5699 = 8'h43 == _t_T_42[31:24] ? 8'h1a : _GEN_5698; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5700 = 8'h44 == _t_T_42[31:24] ? 8'h1b : _GEN_5699; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5701 = 8'h45 == _t_T_42[31:24] ? 8'h6e : _GEN_5700; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5702 = 8'h46 == _t_T_42[31:24] ? 8'h5a : _GEN_5701; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5703 = 8'h47 == _t_T_42[31:24] ? 8'ha0 : _GEN_5702; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5704 = 8'h48 == _t_T_42[31:24] ? 8'h52 : _GEN_5703; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5705 = 8'h49 == _t_T_42[31:24] ? 8'h3b : _GEN_5704; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5706 = 8'h4a == _t_T_42[31:24] ? 8'hd6 : _GEN_5705; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5707 = 8'h4b == _t_T_42[31:24] ? 8'hb3 : _GEN_5706; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5708 = 8'h4c == _t_T_42[31:24] ? 8'h29 : _GEN_5707; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5709 = 8'h4d == _t_T_42[31:24] ? 8'he3 : _GEN_5708; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5710 = 8'h4e == _t_T_42[31:24] ? 8'h2f : _GEN_5709; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5711 = 8'h4f == _t_T_42[31:24] ? 8'h84 : _GEN_5710; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5712 = 8'h50 == _t_T_42[31:24] ? 8'h53 : _GEN_5711; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5713 = 8'h51 == _t_T_42[31:24] ? 8'hd1 : _GEN_5712; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5714 = 8'h52 == _t_T_42[31:24] ? 8'h0 : _GEN_5713; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5715 = 8'h53 == _t_T_42[31:24] ? 8'hed : _GEN_5714; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5716 = 8'h54 == _t_T_42[31:24] ? 8'h20 : _GEN_5715; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5717 = 8'h55 == _t_T_42[31:24] ? 8'hfc : _GEN_5716; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5718 = 8'h56 == _t_T_42[31:24] ? 8'hb1 : _GEN_5717; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5719 = 8'h57 == _t_T_42[31:24] ? 8'h5b : _GEN_5718; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5720 = 8'h58 == _t_T_42[31:24] ? 8'h6a : _GEN_5719; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5721 = 8'h59 == _t_T_42[31:24] ? 8'hcb : _GEN_5720; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5722 = 8'h5a == _t_T_42[31:24] ? 8'hbe : _GEN_5721; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5723 = 8'h5b == _t_T_42[31:24] ? 8'h39 : _GEN_5722; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5724 = 8'h5c == _t_T_42[31:24] ? 8'h4a : _GEN_5723; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5725 = 8'h5d == _t_T_42[31:24] ? 8'h4c : _GEN_5724; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5726 = 8'h5e == _t_T_42[31:24] ? 8'h58 : _GEN_5725; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5727 = 8'h5f == _t_T_42[31:24] ? 8'hcf : _GEN_5726; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5728 = 8'h60 == _t_T_42[31:24] ? 8'hd0 : _GEN_5727; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5729 = 8'h61 == _t_T_42[31:24] ? 8'hef : _GEN_5728; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5730 = 8'h62 == _t_T_42[31:24] ? 8'haa : _GEN_5729; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5731 = 8'h63 == _t_T_42[31:24] ? 8'hfb : _GEN_5730; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5732 = 8'h64 == _t_T_42[31:24] ? 8'h43 : _GEN_5731; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5733 = 8'h65 == _t_T_42[31:24] ? 8'h4d : _GEN_5732; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5734 = 8'h66 == _t_T_42[31:24] ? 8'h33 : _GEN_5733; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5735 = 8'h67 == _t_T_42[31:24] ? 8'h85 : _GEN_5734; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5736 = 8'h68 == _t_T_42[31:24] ? 8'h45 : _GEN_5735; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5737 = 8'h69 == _t_T_42[31:24] ? 8'hf9 : _GEN_5736; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5738 = 8'h6a == _t_T_42[31:24] ? 8'h2 : _GEN_5737; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5739 = 8'h6b == _t_T_42[31:24] ? 8'h7f : _GEN_5738; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5740 = 8'h6c == _t_T_42[31:24] ? 8'h50 : _GEN_5739; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5741 = 8'h6d == _t_T_42[31:24] ? 8'h3c : _GEN_5740; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5742 = 8'h6e == _t_T_42[31:24] ? 8'h9f : _GEN_5741; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5743 = 8'h6f == _t_T_42[31:24] ? 8'ha8 : _GEN_5742; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5744 = 8'h70 == _t_T_42[31:24] ? 8'h51 : _GEN_5743; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5745 = 8'h71 == _t_T_42[31:24] ? 8'ha3 : _GEN_5744; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5746 = 8'h72 == _t_T_42[31:24] ? 8'h40 : _GEN_5745; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5747 = 8'h73 == _t_T_42[31:24] ? 8'h8f : _GEN_5746; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5748 = 8'h74 == _t_T_42[31:24] ? 8'h92 : _GEN_5747; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5749 = 8'h75 == _t_T_42[31:24] ? 8'h9d : _GEN_5748; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5750 = 8'h76 == _t_T_42[31:24] ? 8'h38 : _GEN_5749; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5751 = 8'h77 == _t_T_42[31:24] ? 8'hf5 : _GEN_5750; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5752 = 8'h78 == _t_T_42[31:24] ? 8'hbc : _GEN_5751; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5753 = 8'h79 == _t_T_42[31:24] ? 8'hb6 : _GEN_5752; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5754 = 8'h7a == _t_T_42[31:24] ? 8'hda : _GEN_5753; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5755 = 8'h7b == _t_T_42[31:24] ? 8'h21 : _GEN_5754; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5756 = 8'h7c == _t_T_42[31:24] ? 8'h10 : _GEN_5755; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5757 = 8'h7d == _t_T_42[31:24] ? 8'hff : _GEN_5756; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5758 = 8'h7e == _t_T_42[31:24] ? 8'hf3 : _GEN_5757; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5759 = 8'h7f == _t_T_42[31:24] ? 8'hd2 : _GEN_5758; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5760 = 8'h80 == _t_T_42[31:24] ? 8'hcd : _GEN_5759; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5761 = 8'h81 == _t_T_42[31:24] ? 8'hc : _GEN_5760; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5762 = 8'h82 == _t_T_42[31:24] ? 8'h13 : _GEN_5761; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5763 = 8'h83 == _t_T_42[31:24] ? 8'hec : _GEN_5762; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5764 = 8'h84 == _t_T_42[31:24] ? 8'h5f : _GEN_5763; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5765 = 8'h85 == _t_T_42[31:24] ? 8'h97 : _GEN_5764; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5766 = 8'h86 == _t_T_42[31:24] ? 8'h44 : _GEN_5765; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5767 = 8'h87 == _t_T_42[31:24] ? 8'h17 : _GEN_5766; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5768 = 8'h88 == _t_T_42[31:24] ? 8'hc4 : _GEN_5767; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5769 = 8'h89 == _t_T_42[31:24] ? 8'ha7 : _GEN_5768; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5770 = 8'h8a == _t_T_42[31:24] ? 8'h7e : _GEN_5769; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5771 = 8'h8b == _t_T_42[31:24] ? 8'h3d : _GEN_5770; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5772 = 8'h8c == _t_T_42[31:24] ? 8'h64 : _GEN_5771; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5773 = 8'h8d == _t_T_42[31:24] ? 8'h5d : _GEN_5772; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5774 = 8'h8e == _t_T_42[31:24] ? 8'h19 : _GEN_5773; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5775 = 8'h8f == _t_T_42[31:24] ? 8'h73 : _GEN_5774; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5776 = 8'h90 == _t_T_42[31:24] ? 8'h60 : _GEN_5775; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5777 = 8'h91 == _t_T_42[31:24] ? 8'h81 : _GEN_5776; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5778 = 8'h92 == _t_T_42[31:24] ? 8'h4f : _GEN_5777; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5779 = 8'h93 == _t_T_42[31:24] ? 8'hdc : _GEN_5778; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5780 = 8'h94 == _t_T_42[31:24] ? 8'h22 : _GEN_5779; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5781 = 8'h95 == _t_T_42[31:24] ? 8'h2a : _GEN_5780; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5782 = 8'h96 == _t_T_42[31:24] ? 8'h90 : _GEN_5781; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5783 = 8'h97 == _t_T_42[31:24] ? 8'h88 : _GEN_5782; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5784 = 8'h98 == _t_T_42[31:24] ? 8'h46 : _GEN_5783; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5785 = 8'h99 == _t_T_42[31:24] ? 8'hee : _GEN_5784; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5786 = 8'h9a == _t_T_42[31:24] ? 8'hb8 : _GEN_5785; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5787 = 8'h9b == _t_T_42[31:24] ? 8'h14 : _GEN_5786; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5788 = 8'h9c == _t_T_42[31:24] ? 8'hde : _GEN_5787; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5789 = 8'h9d == _t_T_42[31:24] ? 8'h5e : _GEN_5788; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5790 = 8'h9e == _t_T_42[31:24] ? 8'hb : _GEN_5789; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5791 = 8'h9f == _t_T_42[31:24] ? 8'hdb : _GEN_5790; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5792 = 8'ha0 == _t_T_42[31:24] ? 8'he0 : _GEN_5791; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5793 = 8'ha1 == _t_T_42[31:24] ? 8'h32 : _GEN_5792; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5794 = 8'ha2 == _t_T_42[31:24] ? 8'h3a : _GEN_5793; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5795 = 8'ha3 == _t_T_42[31:24] ? 8'ha : _GEN_5794; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5796 = 8'ha4 == _t_T_42[31:24] ? 8'h49 : _GEN_5795; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5797 = 8'ha5 == _t_T_42[31:24] ? 8'h6 : _GEN_5796; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5798 = 8'ha6 == _t_T_42[31:24] ? 8'h24 : _GEN_5797; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5799 = 8'ha7 == _t_T_42[31:24] ? 8'h5c : _GEN_5798; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5800 = 8'ha8 == _t_T_42[31:24] ? 8'hc2 : _GEN_5799; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5801 = 8'ha9 == _t_T_42[31:24] ? 8'hd3 : _GEN_5800; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5802 = 8'haa == _t_T_42[31:24] ? 8'hac : _GEN_5801; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5803 = 8'hab == _t_T_42[31:24] ? 8'h62 : _GEN_5802; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5804 = 8'hac == _t_T_42[31:24] ? 8'h91 : _GEN_5803; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5805 = 8'had == _t_T_42[31:24] ? 8'h95 : _GEN_5804; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5806 = 8'hae == _t_T_42[31:24] ? 8'he4 : _GEN_5805; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5807 = 8'haf == _t_T_42[31:24] ? 8'h79 : _GEN_5806; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5808 = 8'hb0 == _t_T_42[31:24] ? 8'he7 : _GEN_5807; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5809 = 8'hb1 == _t_T_42[31:24] ? 8'hc8 : _GEN_5808; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5810 = 8'hb2 == _t_T_42[31:24] ? 8'h37 : _GEN_5809; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5811 = 8'hb3 == _t_T_42[31:24] ? 8'h6d : _GEN_5810; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5812 = 8'hb4 == _t_T_42[31:24] ? 8'h8d : _GEN_5811; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5813 = 8'hb5 == _t_T_42[31:24] ? 8'hd5 : _GEN_5812; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5814 = 8'hb6 == _t_T_42[31:24] ? 8'h4e : _GEN_5813; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5815 = 8'hb7 == _t_T_42[31:24] ? 8'ha9 : _GEN_5814; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5816 = 8'hb8 == _t_T_42[31:24] ? 8'h6c : _GEN_5815; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5817 = 8'hb9 == _t_T_42[31:24] ? 8'h56 : _GEN_5816; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5818 = 8'hba == _t_T_42[31:24] ? 8'hf4 : _GEN_5817; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5819 = 8'hbb == _t_T_42[31:24] ? 8'hea : _GEN_5818; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5820 = 8'hbc == _t_T_42[31:24] ? 8'h65 : _GEN_5819; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5821 = 8'hbd == _t_T_42[31:24] ? 8'h7a : _GEN_5820; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5822 = 8'hbe == _t_T_42[31:24] ? 8'hae : _GEN_5821; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5823 = 8'hbf == _t_T_42[31:24] ? 8'h8 : _GEN_5822; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5824 = 8'hc0 == _t_T_42[31:24] ? 8'hba : _GEN_5823; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5825 = 8'hc1 == _t_T_42[31:24] ? 8'h78 : _GEN_5824; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5826 = 8'hc2 == _t_T_42[31:24] ? 8'h25 : _GEN_5825; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5827 = 8'hc3 == _t_T_42[31:24] ? 8'h2e : _GEN_5826; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5828 = 8'hc4 == _t_T_42[31:24] ? 8'h1c : _GEN_5827; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5829 = 8'hc5 == _t_T_42[31:24] ? 8'ha6 : _GEN_5828; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5830 = 8'hc6 == _t_T_42[31:24] ? 8'hb4 : _GEN_5829; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5831 = 8'hc7 == _t_T_42[31:24] ? 8'hc6 : _GEN_5830; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5832 = 8'hc8 == _t_T_42[31:24] ? 8'he8 : _GEN_5831; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5833 = 8'hc9 == _t_T_42[31:24] ? 8'hdd : _GEN_5832; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5834 = 8'hca == _t_T_42[31:24] ? 8'h74 : _GEN_5833; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5835 = 8'hcb == _t_T_42[31:24] ? 8'h1f : _GEN_5834; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5836 = 8'hcc == _t_T_42[31:24] ? 8'h4b : _GEN_5835; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5837 = 8'hcd == _t_T_42[31:24] ? 8'hbd : _GEN_5836; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5838 = 8'hce == _t_T_42[31:24] ? 8'h8b : _GEN_5837; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5839 = 8'hcf == _t_T_42[31:24] ? 8'h8a : _GEN_5838; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5840 = 8'hd0 == _t_T_42[31:24] ? 8'h70 : _GEN_5839; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5841 = 8'hd1 == _t_T_42[31:24] ? 8'h3e : _GEN_5840; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5842 = 8'hd2 == _t_T_42[31:24] ? 8'hb5 : _GEN_5841; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5843 = 8'hd3 == _t_T_42[31:24] ? 8'h66 : _GEN_5842; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5844 = 8'hd4 == _t_T_42[31:24] ? 8'h48 : _GEN_5843; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5845 = 8'hd5 == _t_T_42[31:24] ? 8'h3 : _GEN_5844; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5846 = 8'hd6 == _t_T_42[31:24] ? 8'hf6 : _GEN_5845; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5847 = 8'hd7 == _t_T_42[31:24] ? 8'he : _GEN_5846; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5848 = 8'hd8 == _t_T_42[31:24] ? 8'h61 : _GEN_5847; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5849 = 8'hd9 == _t_T_42[31:24] ? 8'h35 : _GEN_5848; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5850 = 8'hda == _t_T_42[31:24] ? 8'h57 : _GEN_5849; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5851 = 8'hdb == _t_T_42[31:24] ? 8'hb9 : _GEN_5850; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5852 = 8'hdc == _t_T_42[31:24] ? 8'h86 : _GEN_5851; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5853 = 8'hdd == _t_T_42[31:24] ? 8'hc1 : _GEN_5852; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5854 = 8'hde == _t_T_42[31:24] ? 8'h1d : _GEN_5853; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5855 = 8'hdf == _t_T_42[31:24] ? 8'h9e : _GEN_5854; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5856 = 8'he0 == _t_T_42[31:24] ? 8'he1 : _GEN_5855; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5857 = 8'he1 == _t_T_42[31:24] ? 8'hf8 : _GEN_5856; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5858 = 8'he2 == _t_T_42[31:24] ? 8'h98 : _GEN_5857; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5859 = 8'he3 == _t_T_42[31:24] ? 8'h11 : _GEN_5858; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5860 = 8'he4 == _t_T_42[31:24] ? 8'h69 : _GEN_5859; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5861 = 8'he5 == _t_T_42[31:24] ? 8'hd9 : _GEN_5860; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5862 = 8'he6 == _t_T_42[31:24] ? 8'h8e : _GEN_5861; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5863 = 8'he7 == _t_T_42[31:24] ? 8'h94 : _GEN_5862; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5864 = 8'he8 == _t_T_42[31:24] ? 8'h9b : _GEN_5863; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5865 = 8'he9 == _t_T_42[31:24] ? 8'h1e : _GEN_5864; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5866 = 8'hea == _t_T_42[31:24] ? 8'h87 : _GEN_5865; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5867 = 8'heb == _t_T_42[31:24] ? 8'he9 : _GEN_5866; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5868 = 8'hec == _t_T_42[31:24] ? 8'hce : _GEN_5867; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5869 = 8'hed == _t_T_42[31:24] ? 8'h55 : _GEN_5868; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5870 = 8'hee == _t_T_42[31:24] ? 8'h28 : _GEN_5869; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5871 = 8'hef == _t_T_42[31:24] ? 8'hdf : _GEN_5870; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5872 = 8'hf0 == _t_T_42[31:24] ? 8'h8c : _GEN_5871; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5873 = 8'hf1 == _t_T_42[31:24] ? 8'ha1 : _GEN_5872; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5874 = 8'hf2 == _t_T_42[31:24] ? 8'h89 : _GEN_5873; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5875 = 8'hf3 == _t_T_42[31:24] ? 8'hd : _GEN_5874; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5876 = 8'hf4 == _t_T_42[31:24] ? 8'hbf : _GEN_5875; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5877 = 8'hf5 == _t_T_42[31:24] ? 8'he6 : _GEN_5876; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5878 = 8'hf6 == _t_T_42[31:24] ? 8'h42 : _GEN_5877; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5879 = 8'hf7 == _t_T_42[31:24] ? 8'h68 : _GEN_5878; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5880 = 8'hf8 == _t_T_42[31:24] ? 8'h41 : _GEN_5879; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5881 = 8'hf9 == _t_T_42[31:24] ? 8'h99 : _GEN_5880; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5882 = 8'hfa == _t_T_42[31:24] ? 8'h2d : _GEN_5881; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5883 = 8'hfb == _t_T_42[31:24] ? 8'hf : _GEN_5882; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5884 = 8'hfc == _t_T_42[31:24] ? 8'hb0 : _GEN_5883; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5885 = 8'hfd == _t_T_42[31:24] ? 8'h54 : _GEN_5884; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5886 = 8'hfe == _t_T_42[31:24] ? 8'hbb : _GEN_5885; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5887 = 8'hff == _t_T_42[31:24] ? 8'h16 : _GEN_5886; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5889 = 8'h1 == _t_T_42[23:16] ? 8'h7c : 8'h63; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5890 = 8'h2 == _t_T_42[23:16] ? 8'h77 : _GEN_5889; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5891 = 8'h3 == _t_T_42[23:16] ? 8'h7b : _GEN_5890; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5892 = 8'h4 == _t_T_42[23:16] ? 8'hf2 : _GEN_5891; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5893 = 8'h5 == _t_T_42[23:16] ? 8'h6b : _GEN_5892; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5894 = 8'h6 == _t_T_42[23:16] ? 8'h6f : _GEN_5893; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5895 = 8'h7 == _t_T_42[23:16] ? 8'hc5 : _GEN_5894; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5896 = 8'h8 == _t_T_42[23:16] ? 8'h30 : _GEN_5895; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5897 = 8'h9 == _t_T_42[23:16] ? 8'h1 : _GEN_5896; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5898 = 8'ha == _t_T_42[23:16] ? 8'h67 : _GEN_5897; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5899 = 8'hb == _t_T_42[23:16] ? 8'h2b : _GEN_5898; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5900 = 8'hc == _t_T_42[23:16] ? 8'hfe : _GEN_5899; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5901 = 8'hd == _t_T_42[23:16] ? 8'hd7 : _GEN_5900; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5902 = 8'he == _t_T_42[23:16] ? 8'hab : _GEN_5901; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5903 = 8'hf == _t_T_42[23:16] ? 8'h76 : _GEN_5902; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5904 = 8'h10 == _t_T_42[23:16] ? 8'hca : _GEN_5903; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5905 = 8'h11 == _t_T_42[23:16] ? 8'h82 : _GEN_5904; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5906 = 8'h12 == _t_T_42[23:16] ? 8'hc9 : _GEN_5905; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5907 = 8'h13 == _t_T_42[23:16] ? 8'h7d : _GEN_5906; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5908 = 8'h14 == _t_T_42[23:16] ? 8'hfa : _GEN_5907; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5909 = 8'h15 == _t_T_42[23:16] ? 8'h59 : _GEN_5908; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5910 = 8'h16 == _t_T_42[23:16] ? 8'h47 : _GEN_5909; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5911 = 8'h17 == _t_T_42[23:16] ? 8'hf0 : _GEN_5910; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5912 = 8'h18 == _t_T_42[23:16] ? 8'had : _GEN_5911; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5913 = 8'h19 == _t_T_42[23:16] ? 8'hd4 : _GEN_5912; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5914 = 8'h1a == _t_T_42[23:16] ? 8'ha2 : _GEN_5913; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5915 = 8'h1b == _t_T_42[23:16] ? 8'haf : _GEN_5914; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5916 = 8'h1c == _t_T_42[23:16] ? 8'h9c : _GEN_5915; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5917 = 8'h1d == _t_T_42[23:16] ? 8'ha4 : _GEN_5916; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5918 = 8'h1e == _t_T_42[23:16] ? 8'h72 : _GEN_5917; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5919 = 8'h1f == _t_T_42[23:16] ? 8'hc0 : _GEN_5918; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5920 = 8'h20 == _t_T_42[23:16] ? 8'hb7 : _GEN_5919; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5921 = 8'h21 == _t_T_42[23:16] ? 8'hfd : _GEN_5920; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5922 = 8'h22 == _t_T_42[23:16] ? 8'h93 : _GEN_5921; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5923 = 8'h23 == _t_T_42[23:16] ? 8'h26 : _GEN_5922; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5924 = 8'h24 == _t_T_42[23:16] ? 8'h36 : _GEN_5923; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5925 = 8'h25 == _t_T_42[23:16] ? 8'h3f : _GEN_5924; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5926 = 8'h26 == _t_T_42[23:16] ? 8'hf7 : _GEN_5925; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5927 = 8'h27 == _t_T_42[23:16] ? 8'hcc : _GEN_5926; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5928 = 8'h28 == _t_T_42[23:16] ? 8'h34 : _GEN_5927; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5929 = 8'h29 == _t_T_42[23:16] ? 8'ha5 : _GEN_5928; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5930 = 8'h2a == _t_T_42[23:16] ? 8'he5 : _GEN_5929; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5931 = 8'h2b == _t_T_42[23:16] ? 8'hf1 : _GEN_5930; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5932 = 8'h2c == _t_T_42[23:16] ? 8'h71 : _GEN_5931; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5933 = 8'h2d == _t_T_42[23:16] ? 8'hd8 : _GEN_5932; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5934 = 8'h2e == _t_T_42[23:16] ? 8'h31 : _GEN_5933; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5935 = 8'h2f == _t_T_42[23:16] ? 8'h15 : _GEN_5934; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5936 = 8'h30 == _t_T_42[23:16] ? 8'h4 : _GEN_5935; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5937 = 8'h31 == _t_T_42[23:16] ? 8'hc7 : _GEN_5936; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5938 = 8'h32 == _t_T_42[23:16] ? 8'h23 : _GEN_5937; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5939 = 8'h33 == _t_T_42[23:16] ? 8'hc3 : _GEN_5938; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5940 = 8'h34 == _t_T_42[23:16] ? 8'h18 : _GEN_5939; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5941 = 8'h35 == _t_T_42[23:16] ? 8'h96 : _GEN_5940; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5942 = 8'h36 == _t_T_42[23:16] ? 8'h5 : _GEN_5941; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5943 = 8'h37 == _t_T_42[23:16] ? 8'h9a : _GEN_5942; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5944 = 8'h38 == _t_T_42[23:16] ? 8'h7 : _GEN_5943; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5945 = 8'h39 == _t_T_42[23:16] ? 8'h12 : _GEN_5944; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5946 = 8'h3a == _t_T_42[23:16] ? 8'h80 : _GEN_5945; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5947 = 8'h3b == _t_T_42[23:16] ? 8'he2 : _GEN_5946; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5948 = 8'h3c == _t_T_42[23:16] ? 8'heb : _GEN_5947; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5949 = 8'h3d == _t_T_42[23:16] ? 8'h27 : _GEN_5948; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5950 = 8'h3e == _t_T_42[23:16] ? 8'hb2 : _GEN_5949; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5951 = 8'h3f == _t_T_42[23:16] ? 8'h75 : _GEN_5950; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5952 = 8'h40 == _t_T_42[23:16] ? 8'h9 : _GEN_5951; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5953 = 8'h41 == _t_T_42[23:16] ? 8'h83 : _GEN_5952; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5954 = 8'h42 == _t_T_42[23:16] ? 8'h2c : _GEN_5953; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5955 = 8'h43 == _t_T_42[23:16] ? 8'h1a : _GEN_5954; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5956 = 8'h44 == _t_T_42[23:16] ? 8'h1b : _GEN_5955; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5957 = 8'h45 == _t_T_42[23:16] ? 8'h6e : _GEN_5956; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5958 = 8'h46 == _t_T_42[23:16] ? 8'h5a : _GEN_5957; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5959 = 8'h47 == _t_T_42[23:16] ? 8'ha0 : _GEN_5958; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5960 = 8'h48 == _t_T_42[23:16] ? 8'h52 : _GEN_5959; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5961 = 8'h49 == _t_T_42[23:16] ? 8'h3b : _GEN_5960; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5962 = 8'h4a == _t_T_42[23:16] ? 8'hd6 : _GEN_5961; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5963 = 8'h4b == _t_T_42[23:16] ? 8'hb3 : _GEN_5962; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5964 = 8'h4c == _t_T_42[23:16] ? 8'h29 : _GEN_5963; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5965 = 8'h4d == _t_T_42[23:16] ? 8'he3 : _GEN_5964; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5966 = 8'h4e == _t_T_42[23:16] ? 8'h2f : _GEN_5965; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5967 = 8'h4f == _t_T_42[23:16] ? 8'h84 : _GEN_5966; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5968 = 8'h50 == _t_T_42[23:16] ? 8'h53 : _GEN_5967; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5969 = 8'h51 == _t_T_42[23:16] ? 8'hd1 : _GEN_5968; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5970 = 8'h52 == _t_T_42[23:16] ? 8'h0 : _GEN_5969; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5971 = 8'h53 == _t_T_42[23:16] ? 8'hed : _GEN_5970; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5972 = 8'h54 == _t_T_42[23:16] ? 8'h20 : _GEN_5971; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5973 = 8'h55 == _t_T_42[23:16] ? 8'hfc : _GEN_5972; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5974 = 8'h56 == _t_T_42[23:16] ? 8'hb1 : _GEN_5973; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5975 = 8'h57 == _t_T_42[23:16] ? 8'h5b : _GEN_5974; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5976 = 8'h58 == _t_T_42[23:16] ? 8'h6a : _GEN_5975; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5977 = 8'h59 == _t_T_42[23:16] ? 8'hcb : _GEN_5976; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5978 = 8'h5a == _t_T_42[23:16] ? 8'hbe : _GEN_5977; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5979 = 8'h5b == _t_T_42[23:16] ? 8'h39 : _GEN_5978; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5980 = 8'h5c == _t_T_42[23:16] ? 8'h4a : _GEN_5979; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5981 = 8'h5d == _t_T_42[23:16] ? 8'h4c : _GEN_5980; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5982 = 8'h5e == _t_T_42[23:16] ? 8'h58 : _GEN_5981; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5983 = 8'h5f == _t_T_42[23:16] ? 8'hcf : _GEN_5982; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5984 = 8'h60 == _t_T_42[23:16] ? 8'hd0 : _GEN_5983; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5985 = 8'h61 == _t_T_42[23:16] ? 8'hef : _GEN_5984; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5986 = 8'h62 == _t_T_42[23:16] ? 8'haa : _GEN_5985; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5987 = 8'h63 == _t_T_42[23:16] ? 8'hfb : _GEN_5986; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5988 = 8'h64 == _t_T_42[23:16] ? 8'h43 : _GEN_5987; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5989 = 8'h65 == _t_T_42[23:16] ? 8'h4d : _GEN_5988; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5990 = 8'h66 == _t_T_42[23:16] ? 8'h33 : _GEN_5989; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5991 = 8'h67 == _t_T_42[23:16] ? 8'h85 : _GEN_5990; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5992 = 8'h68 == _t_T_42[23:16] ? 8'h45 : _GEN_5991; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5993 = 8'h69 == _t_T_42[23:16] ? 8'hf9 : _GEN_5992; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5994 = 8'h6a == _t_T_42[23:16] ? 8'h2 : _GEN_5993; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5995 = 8'h6b == _t_T_42[23:16] ? 8'h7f : _GEN_5994; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5996 = 8'h6c == _t_T_42[23:16] ? 8'h50 : _GEN_5995; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5997 = 8'h6d == _t_T_42[23:16] ? 8'h3c : _GEN_5996; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5998 = 8'h6e == _t_T_42[23:16] ? 8'h9f : _GEN_5997; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_5999 = 8'h6f == _t_T_42[23:16] ? 8'ha8 : _GEN_5998; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6000 = 8'h70 == _t_T_42[23:16] ? 8'h51 : _GEN_5999; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6001 = 8'h71 == _t_T_42[23:16] ? 8'ha3 : _GEN_6000; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6002 = 8'h72 == _t_T_42[23:16] ? 8'h40 : _GEN_6001; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6003 = 8'h73 == _t_T_42[23:16] ? 8'h8f : _GEN_6002; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6004 = 8'h74 == _t_T_42[23:16] ? 8'h92 : _GEN_6003; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6005 = 8'h75 == _t_T_42[23:16] ? 8'h9d : _GEN_6004; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6006 = 8'h76 == _t_T_42[23:16] ? 8'h38 : _GEN_6005; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6007 = 8'h77 == _t_T_42[23:16] ? 8'hf5 : _GEN_6006; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6008 = 8'h78 == _t_T_42[23:16] ? 8'hbc : _GEN_6007; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6009 = 8'h79 == _t_T_42[23:16] ? 8'hb6 : _GEN_6008; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6010 = 8'h7a == _t_T_42[23:16] ? 8'hda : _GEN_6009; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6011 = 8'h7b == _t_T_42[23:16] ? 8'h21 : _GEN_6010; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6012 = 8'h7c == _t_T_42[23:16] ? 8'h10 : _GEN_6011; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6013 = 8'h7d == _t_T_42[23:16] ? 8'hff : _GEN_6012; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6014 = 8'h7e == _t_T_42[23:16] ? 8'hf3 : _GEN_6013; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6015 = 8'h7f == _t_T_42[23:16] ? 8'hd2 : _GEN_6014; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6016 = 8'h80 == _t_T_42[23:16] ? 8'hcd : _GEN_6015; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6017 = 8'h81 == _t_T_42[23:16] ? 8'hc : _GEN_6016; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6018 = 8'h82 == _t_T_42[23:16] ? 8'h13 : _GEN_6017; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6019 = 8'h83 == _t_T_42[23:16] ? 8'hec : _GEN_6018; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6020 = 8'h84 == _t_T_42[23:16] ? 8'h5f : _GEN_6019; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6021 = 8'h85 == _t_T_42[23:16] ? 8'h97 : _GEN_6020; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6022 = 8'h86 == _t_T_42[23:16] ? 8'h44 : _GEN_6021; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6023 = 8'h87 == _t_T_42[23:16] ? 8'h17 : _GEN_6022; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6024 = 8'h88 == _t_T_42[23:16] ? 8'hc4 : _GEN_6023; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6025 = 8'h89 == _t_T_42[23:16] ? 8'ha7 : _GEN_6024; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6026 = 8'h8a == _t_T_42[23:16] ? 8'h7e : _GEN_6025; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6027 = 8'h8b == _t_T_42[23:16] ? 8'h3d : _GEN_6026; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6028 = 8'h8c == _t_T_42[23:16] ? 8'h64 : _GEN_6027; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6029 = 8'h8d == _t_T_42[23:16] ? 8'h5d : _GEN_6028; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6030 = 8'h8e == _t_T_42[23:16] ? 8'h19 : _GEN_6029; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6031 = 8'h8f == _t_T_42[23:16] ? 8'h73 : _GEN_6030; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6032 = 8'h90 == _t_T_42[23:16] ? 8'h60 : _GEN_6031; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6033 = 8'h91 == _t_T_42[23:16] ? 8'h81 : _GEN_6032; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6034 = 8'h92 == _t_T_42[23:16] ? 8'h4f : _GEN_6033; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6035 = 8'h93 == _t_T_42[23:16] ? 8'hdc : _GEN_6034; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6036 = 8'h94 == _t_T_42[23:16] ? 8'h22 : _GEN_6035; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6037 = 8'h95 == _t_T_42[23:16] ? 8'h2a : _GEN_6036; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6038 = 8'h96 == _t_T_42[23:16] ? 8'h90 : _GEN_6037; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6039 = 8'h97 == _t_T_42[23:16] ? 8'h88 : _GEN_6038; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6040 = 8'h98 == _t_T_42[23:16] ? 8'h46 : _GEN_6039; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6041 = 8'h99 == _t_T_42[23:16] ? 8'hee : _GEN_6040; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6042 = 8'h9a == _t_T_42[23:16] ? 8'hb8 : _GEN_6041; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6043 = 8'h9b == _t_T_42[23:16] ? 8'h14 : _GEN_6042; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6044 = 8'h9c == _t_T_42[23:16] ? 8'hde : _GEN_6043; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6045 = 8'h9d == _t_T_42[23:16] ? 8'h5e : _GEN_6044; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6046 = 8'h9e == _t_T_42[23:16] ? 8'hb : _GEN_6045; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6047 = 8'h9f == _t_T_42[23:16] ? 8'hdb : _GEN_6046; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6048 = 8'ha0 == _t_T_42[23:16] ? 8'he0 : _GEN_6047; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6049 = 8'ha1 == _t_T_42[23:16] ? 8'h32 : _GEN_6048; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6050 = 8'ha2 == _t_T_42[23:16] ? 8'h3a : _GEN_6049; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6051 = 8'ha3 == _t_T_42[23:16] ? 8'ha : _GEN_6050; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6052 = 8'ha4 == _t_T_42[23:16] ? 8'h49 : _GEN_6051; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6053 = 8'ha5 == _t_T_42[23:16] ? 8'h6 : _GEN_6052; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6054 = 8'ha6 == _t_T_42[23:16] ? 8'h24 : _GEN_6053; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6055 = 8'ha7 == _t_T_42[23:16] ? 8'h5c : _GEN_6054; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6056 = 8'ha8 == _t_T_42[23:16] ? 8'hc2 : _GEN_6055; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6057 = 8'ha9 == _t_T_42[23:16] ? 8'hd3 : _GEN_6056; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6058 = 8'haa == _t_T_42[23:16] ? 8'hac : _GEN_6057; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6059 = 8'hab == _t_T_42[23:16] ? 8'h62 : _GEN_6058; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6060 = 8'hac == _t_T_42[23:16] ? 8'h91 : _GEN_6059; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6061 = 8'had == _t_T_42[23:16] ? 8'h95 : _GEN_6060; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6062 = 8'hae == _t_T_42[23:16] ? 8'he4 : _GEN_6061; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6063 = 8'haf == _t_T_42[23:16] ? 8'h79 : _GEN_6062; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6064 = 8'hb0 == _t_T_42[23:16] ? 8'he7 : _GEN_6063; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6065 = 8'hb1 == _t_T_42[23:16] ? 8'hc8 : _GEN_6064; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6066 = 8'hb2 == _t_T_42[23:16] ? 8'h37 : _GEN_6065; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6067 = 8'hb3 == _t_T_42[23:16] ? 8'h6d : _GEN_6066; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6068 = 8'hb4 == _t_T_42[23:16] ? 8'h8d : _GEN_6067; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6069 = 8'hb5 == _t_T_42[23:16] ? 8'hd5 : _GEN_6068; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6070 = 8'hb6 == _t_T_42[23:16] ? 8'h4e : _GEN_6069; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6071 = 8'hb7 == _t_T_42[23:16] ? 8'ha9 : _GEN_6070; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6072 = 8'hb8 == _t_T_42[23:16] ? 8'h6c : _GEN_6071; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6073 = 8'hb9 == _t_T_42[23:16] ? 8'h56 : _GEN_6072; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6074 = 8'hba == _t_T_42[23:16] ? 8'hf4 : _GEN_6073; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6075 = 8'hbb == _t_T_42[23:16] ? 8'hea : _GEN_6074; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6076 = 8'hbc == _t_T_42[23:16] ? 8'h65 : _GEN_6075; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6077 = 8'hbd == _t_T_42[23:16] ? 8'h7a : _GEN_6076; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6078 = 8'hbe == _t_T_42[23:16] ? 8'hae : _GEN_6077; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6079 = 8'hbf == _t_T_42[23:16] ? 8'h8 : _GEN_6078; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6080 = 8'hc0 == _t_T_42[23:16] ? 8'hba : _GEN_6079; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6081 = 8'hc1 == _t_T_42[23:16] ? 8'h78 : _GEN_6080; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6082 = 8'hc2 == _t_T_42[23:16] ? 8'h25 : _GEN_6081; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6083 = 8'hc3 == _t_T_42[23:16] ? 8'h2e : _GEN_6082; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6084 = 8'hc4 == _t_T_42[23:16] ? 8'h1c : _GEN_6083; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6085 = 8'hc5 == _t_T_42[23:16] ? 8'ha6 : _GEN_6084; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6086 = 8'hc6 == _t_T_42[23:16] ? 8'hb4 : _GEN_6085; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6087 = 8'hc7 == _t_T_42[23:16] ? 8'hc6 : _GEN_6086; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6088 = 8'hc8 == _t_T_42[23:16] ? 8'he8 : _GEN_6087; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6089 = 8'hc9 == _t_T_42[23:16] ? 8'hdd : _GEN_6088; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6090 = 8'hca == _t_T_42[23:16] ? 8'h74 : _GEN_6089; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6091 = 8'hcb == _t_T_42[23:16] ? 8'h1f : _GEN_6090; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6092 = 8'hcc == _t_T_42[23:16] ? 8'h4b : _GEN_6091; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6093 = 8'hcd == _t_T_42[23:16] ? 8'hbd : _GEN_6092; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6094 = 8'hce == _t_T_42[23:16] ? 8'h8b : _GEN_6093; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6095 = 8'hcf == _t_T_42[23:16] ? 8'h8a : _GEN_6094; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6096 = 8'hd0 == _t_T_42[23:16] ? 8'h70 : _GEN_6095; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6097 = 8'hd1 == _t_T_42[23:16] ? 8'h3e : _GEN_6096; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6098 = 8'hd2 == _t_T_42[23:16] ? 8'hb5 : _GEN_6097; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6099 = 8'hd3 == _t_T_42[23:16] ? 8'h66 : _GEN_6098; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6100 = 8'hd4 == _t_T_42[23:16] ? 8'h48 : _GEN_6099; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6101 = 8'hd5 == _t_T_42[23:16] ? 8'h3 : _GEN_6100; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6102 = 8'hd6 == _t_T_42[23:16] ? 8'hf6 : _GEN_6101; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6103 = 8'hd7 == _t_T_42[23:16] ? 8'he : _GEN_6102; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6104 = 8'hd8 == _t_T_42[23:16] ? 8'h61 : _GEN_6103; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6105 = 8'hd9 == _t_T_42[23:16] ? 8'h35 : _GEN_6104; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6106 = 8'hda == _t_T_42[23:16] ? 8'h57 : _GEN_6105; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6107 = 8'hdb == _t_T_42[23:16] ? 8'hb9 : _GEN_6106; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6108 = 8'hdc == _t_T_42[23:16] ? 8'h86 : _GEN_6107; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6109 = 8'hdd == _t_T_42[23:16] ? 8'hc1 : _GEN_6108; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6110 = 8'hde == _t_T_42[23:16] ? 8'h1d : _GEN_6109; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6111 = 8'hdf == _t_T_42[23:16] ? 8'h9e : _GEN_6110; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6112 = 8'he0 == _t_T_42[23:16] ? 8'he1 : _GEN_6111; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6113 = 8'he1 == _t_T_42[23:16] ? 8'hf8 : _GEN_6112; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6114 = 8'he2 == _t_T_42[23:16] ? 8'h98 : _GEN_6113; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6115 = 8'he3 == _t_T_42[23:16] ? 8'h11 : _GEN_6114; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6116 = 8'he4 == _t_T_42[23:16] ? 8'h69 : _GEN_6115; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6117 = 8'he5 == _t_T_42[23:16] ? 8'hd9 : _GEN_6116; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6118 = 8'he6 == _t_T_42[23:16] ? 8'h8e : _GEN_6117; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6119 = 8'he7 == _t_T_42[23:16] ? 8'h94 : _GEN_6118; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6120 = 8'he8 == _t_T_42[23:16] ? 8'h9b : _GEN_6119; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6121 = 8'he9 == _t_T_42[23:16] ? 8'h1e : _GEN_6120; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6122 = 8'hea == _t_T_42[23:16] ? 8'h87 : _GEN_6121; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6123 = 8'heb == _t_T_42[23:16] ? 8'he9 : _GEN_6122; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6124 = 8'hec == _t_T_42[23:16] ? 8'hce : _GEN_6123; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6125 = 8'hed == _t_T_42[23:16] ? 8'h55 : _GEN_6124; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6126 = 8'hee == _t_T_42[23:16] ? 8'h28 : _GEN_6125; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6127 = 8'hef == _t_T_42[23:16] ? 8'hdf : _GEN_6126; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6128 = 8'hf0 == _t_T_42[23:16] ? 8'h8c : _GEN_6127; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6129 = 8'hf1 == _t_T_42[23:16] ? 8'ha1 : _GEN_6128; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6130 = 8'hf2 == _t_T_42[23:16] ? 8'h89 : _GEN_6129; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6131 = 8'hf3 == _t_T_42[23:16] ? 8'hd : _GEN_6130; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6132 = 8'hf4 == _t_T_42[23:16] ? 8'hbf : _GEN_6131; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6133 = 8'hf5 == _t_T_42[23:16] ? 8'he6 : _GEN_6132; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6134 = 8'hf6 == _t_T_42[23:16] ? 8'h42 : _GEN_6133; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6135 = 8'hf7 == _t_T_42[23:16] ? 8'h68 : _GEN_6134; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6136 = 8'hf8 == _t_T_42[23:16] ? 8'h41 : _GEN_6135; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6137 = 8'hf9 == _t_T_42[23:16] ? 8'h99 : _GEN_6136; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6138 = 8'hfa == _t_T_42[23:16] ? 8'h2d : _GEN_6137; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6139 = 8'hfb == _t_T_42[23:16] ? 8'hf : _GEN_6138; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6140 = 8'hfc == _t_T_42[23:16] ? 8'hb0 : _GEN_6139; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6141 = 8'hfd == _t_T_42[23:16] ? 8'h54 : _GEN_6140; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6142 = 8'hfe == _t_T_42[23:16] ? 8'hbb : _GEN_6141; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6143 = 8'hff == _t_T_42[23:16] ? 8'h16 : _GEN_6142; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [31:0] _t_T_47 = {_GEN_5887,_GEN_6143,_GEN_5375,_GEN_5631}; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:8]
  wire [31:0] t_5 = _t_T_47 ^ 32'h20000000; // @[src/main/scala/crypto/aes/KeySchedule.scala 59:32]
  wire [31:0] w_24 = w_20 ^ t_5; // @[src/main/scala/crypto/aes/KeySchedule.scala 63:21]
  wire [31:0] w_25 = w_21 ^ w_24; // @[src/main/scala/crypto/aes/KeySchedule.scala 63:21]
  wire [31:0] w_26 = w_22 ^ w_25; // @[src/main/scala/crypto/aes/KeySchedule.scala 63:21]
  wire [31:0] w_27 = w_23 ^ w_26; // @[src/main/scala/crypto/aes/KeySchedule.scala 63:21]
  wire [31:0] _t_T_50 = {w_27[23:0],w_27[31:24]}; // @[src/main/scala/crypto/aes/KeySchedule.scala 23:43]
  wire [7:0] _GEN_6145 = 8'h1 == _t_T_50[15:8] ? 8'h7c : 8'h63; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6146 = 8'h2 == _t_T_50[15:8] ? 8'h77 : _GEN_6145; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6147 = 8'h3 == _t_T_50[15:8] ? 8'h7b : _GEN_6146; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6148 = 8'h4 == _t_T_50[15:8] ? 8'hf2 : _GEN_6147; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6149 = 8'h5 == _t_T_50[15:8] ? 8'h6b : _GEN_6148; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6150 = 8'h6 == _t_T_50[15:8] ? 8'h6f : _GEN_6149; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6151 = 8'h7 == _t_T_50[15:8] ? 8'hc5 : _GEN_6150; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6152 = 8'h8 == _t_T_50[15:8] ? 8'h30 : _GEN_6151; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6153 = 8'h9 == _t_T_50[15:8] ? 8'h1 : _GEN_6152; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6154 = 8'ha == _t_T_50[15:8] ? 8'h67 : _GEN_6153; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6155 = 8'hb == _t_T_50[15:8] ? 8'h2b : _GEN_6154; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6156 = 8'hc == _t_T_50[15:8] ? 8'hfe : _GEN_6155; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6157 = 8'hd == _t_T_50[15:8] ? 8'hd7 : _GEN_6156; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6158 = 8'he == _t_T_50[15:8] ? 8'hab : _GEN_6157; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6159 = 8'hf == _t_T_50[15:8] ? 8'h76 : _GEN_6158; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6160 = 8'h10 == _t_T_50[15:8] ? 8'hca : _GEN_6159; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6161 = 8'h11 == _t_T_50[15:8] ? 8'h82 : _GEN_6160; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6162 = 8'h12 == _t_T_50[15:8] ? 8'hc9 : _GEN_6161; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6163 = 8'h13 == _t_T_50[15:8] ? 8'h7d : _GEN_6162; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6164 = 8'h14 == _t_T_50[15:8] ? 8'hfa : _GEN_6163; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6165 = 8'h15 == _t_T_50[15:8] ? 8'h59 : _GEN_6164; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6166 = 8'h16 == _t_T_50[15:8] ? 8'h47 : _GEN_6165; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6167 = 8'h17 == _t_T_50[15:8] ? 8'hf0 : _GEN_6166; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6168 = 8'h18 == _t_T_50[15:8] ? 8'had : _GEN_6167; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6169 = 8'h19 == _t_T_50[15:8] ? 8'hd4 : _GEN_6168; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6170 = 8'h1a == _t_T_50[15:8] ? 8'ha2 : _GEN_6169; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6171 = 8'h1b == _t_T_50[15:8] ? 8'haf : _GEN_6170; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6172 = 8'h1c == _t_T_50[15:8] ? 8'h9c : _GEN_6171; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6173 = 8'h1d == _t_T_50[15:8] ? 8'ha4 : _GEN_6172; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6174 = 8'h1e == _t_T_50[15:8] ? 8'h72 : _GEN_6173; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6175 = 8'h1f == _t_T_50[15:8] ? 8'hc0 : _GEN_6174; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6176 = 8'h20 == _t_T_50[15:8] ? 8'hb7 : _GEN_6175; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6177 = 8'h21 == _t_T_50[15:8] ? 8'hfd : _GEN_6176; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6178 = 8'h22 == _t_T_50[15:8] ? 8'h93 : _GEN_6177; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6179 = 8'h23 == _t_T_50[15:8] ? 8'h26 : _GEN_6178; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6180 = 8'h24 == _t_T_50[15:8] ? 8'h36 : _GEN_6179; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6181 = 8'h25 == _t_T_50[15:8] ? 8'h3f : _GEN_6180; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6182 = 8'h26 == _t_T_50[15:8] ? 8'hf7 : _GEN_6181; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6183 = 8'h27 == _t_T_50[15:8] ? 8'hcc : _GEN_6182; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6184 = 8'h28 == _t_T_50[15:8] ? 8'h34 : _GEN_6183; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6185 = 8'h29 == _t_T_50[15:8] ? 8'ha5 : _GEN_6184; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6186 = 8'h2a == _t_T_50[15:8] ? 8'he5 : _GEN_6185; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6187 = 8'h2b == _t_T_50[15:8] ? 8'hf1 : _GEN_6186; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6188 = 8'h2c == _t_T_50[15:8] ? 8'h71 : _GEN_6187; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6189 = 8'h2d == _t_T_50[15:8] ? 8'hd8 : _GEN_6188; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6190 = 8'h2e == _t_T_50[15:8] ? 8'h31 : _GEN_6189; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6191 = 8'h2f == _t_T_50[15:8] ? 8'h15 : _GEN_6190; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6192 = 8'h30 == _t_T_50[15:8] ? 8'h4 : _GEN_6191; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6193 = 8'h31 == _t_T_50[15:8] ? 8'hc7 : _GEN_6192; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6194 = 8'h32 == _t_T_50[15:8] ? 8'h23 : _GEN_6193; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6195 = 8'h33 == _t_T_50[15:8] ? 8'hc3 : _GEN_6194; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6196 = 8'h34 == _t_T_50[15:8] ? 8'h18 : _GEN_6195; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6197 = 8'h35 == _t_T_50[15:8] ? 8'h96 : _GEN_6196; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6198 = 8'h36 == _t_T_50[15:8] ? 8'h5 : _GEN_6197; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6199 = 8'h37 == _t_T_50[15:8] ? 8'h9a : _GEN_6198; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6200 = 8'h38 == _t_T_50[15:8] ? 8'h7 : _GEN_6199; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6201 = 8'h39 == _t_T_50[15:8] ? 8'h12 : _GEN_6200; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6202 = 8'h3a == _t_T_50[15:8] ? 8'h80 : _GEN_6201; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6203 = 8'h3b == _t_T_50[15:8] ? 8'he2 : _GEN_6202; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6204 = 8'h3c == _t_T_50[15:8] ? 8'heb : _GEN_6203; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6205 = 8'h3d == _t_T_50[15:8] ? 8'h27 : _GEN_6204; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6206 = 8'h3e == _t_T_50[15:8] ? 8'hb2 : _GEN_6205; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6207 = 8'h3f == _t_T_50[15:8] ? 8'h75 : _GEN_6206; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6208 = 8'h40 == _t_T_50[15:8] ? 8'h9 : _GEN_6207; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6209 = 8'h41 == _t_T_50[15:8] ? 8'h83 : _GEN_6208; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6210 = 8'h42 == _t_T_50[15:8] ? 8'h2c : _GEN_6209; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6211 = 8'h43 == _t_T_50[15:8] ? 8'h1a : _GEN_6210; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6212 = 8'h44 == _t_T_50[15:8] ? 8'h1b : _GEN_6211; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6213 = 8'h45 == _t_T_50[15:8] ? 8'h6e : _GEN_6212; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6214 = 8'h46 == _t_T_50[15:8] ? 8'h5a : _GEN_6213; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6215 = 8'h47 == _t_T_50[15:8] ? 8'ha0 : _GEN_6214; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6216 = 8'h48 == _t_T_50[15:8] ? 8'h52 : _GEN_6215; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6217 = 8'h49 == _t_T_50[15:8] ? 8'h3b : _GEN_6216; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6218 = 8'h4a == _t_T_50[15:8] ? 8'hd6 : _GEN_6217; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6219 = 8'h4b == _t_T_50[15:8] ? 8'hb3 : _GEN_6218; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6220 = 8'h4c == _t_T_50[15:8] ? 8'h29 : _GEN_6219; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6221 = 8'h4d == _t_T_50[15:8] ? 8'he3 : _GEN_6220; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6222 = 8'h4e == _t_T_50[15:8] ? 8'h2f : _GEN_6221; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6223 = 8'h4f == _t_T_50[15:8] ? 8'h84 : _GEN_6222; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6224 = 8'h50 == _t_T_50[15:8] ? 8'h53 : _GEN_6223; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6225 = 8'h51 == _t_T_50[15:8] ? 8'hd1 : _GEN_6224; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6226 = 8'h52 == _t_T_50[15:8] ? 8'h0 : _GEN_6225; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6227 = 8'h53 == _t_T_50[15:8] ? 8'hed : _GEN_6226; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6228 = 8'h54 == _t_T_50[15:8] ? 8'h20 : _GEN_6227; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6229 = 8'h55 == _t_T_50[15:8] ? 8'hfc : _GEN_6228; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6230 = 8'h56 == _t_T_50[15:8] ? 8'hb1 : _GEN_6229; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6231 = 8'h57 == _t_T_50[15:8] ? 8'h5b : _GEN_6230; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6232 = 8'h58 == _t_T_50[15:8] ? 8'h6a : _GEN_6231; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6233 = 8'h59 == _t_T_50[15:8] ? 8'hcb : _GEN_6232; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6234 = 8'h5a == _t_T_50[15:8] ? 8'hbe : _GEN_6233; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6235 = 8'h5b == _t_T_50[15:8] ? 8'h39 : _GEN_6234; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6236 = 8'h5c == _t_T_50[15:8] ? 8'h4a : _GEN_6235; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6237 = 8'h5d == _t_T_50[15:8] ? 8'h4c : _GEN_6236; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6238 = 8'h5e == _t_T_50[15:8] ? 8'h58 : _GEN_6237; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6239 = 8'h5f == _t_T_50[15:8] ? 8'hcf : _GEN_6238; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6240 = 8'h60 == _t_T_50[15:8] ? 8'hd0 : _GEN_6239; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6241 = 8'h61 == _t_T_50[15:8] ? 8'hef : _GEN_6240; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6242 = 8'h62 == _t_T_50[15:8] ? 8'haa : _GEN_6241; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6243 = 8'h63 == _t_T_50[15:8] ? 8'hfb : _GEN_6242; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6244 = 8'h64 == _t_T_50[15:8] ? 8'h43 : _GEN_6243; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6245 = 8'h65 == _t_T_50[15:8] ? 8'h4d : _GEN_6244; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6246 = 8'h66 == _t_T_50[15:8] ? 8'h33 : _GEN_6245; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6247 = 8'h67 == _t_T_50[15:8] ? 8'h85 : _GEN_6246; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6248 = 8'h68 == _t_T_50[15:8] ? 8'h45 : _GEN_6247; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6249 = 8'h69 == _t_T_50[15:8] ? 8'hf9 : _GEN_6248; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6250 = 8'h6a == _t_T_50[15:8] ? 8'h2 : _GEN_6249; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6251 = 8'h6b == _t_T_50[15:8] ? 8'h7f : _GEN_6250; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6252 = 8'h6c == _t_T_50[15:8] ? 8'h50 : _GEN_6251; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6253 = 8'h6d == _t_T_50[15:8] ? 8'h3c : _GEN_6252; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6254 = 8'h6e == _t_T_50[15:8] ? 8'h9f : _GEN_6253; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6255 = 8'h6f == _t_T_50[15:8] ? 8'ha8 : _GEN_6254; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6256 = 8'h70 == _t_T_50[15:8] ? 8'h51 : _GEN_6255; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6257 = 8'h71 == _t_T_50[15:8] ? 8'ha3 : _GEN_6256; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6258 = 8'h72 == _t_T_50[15:8] ? 8'h40 : _GEN_6257; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6259 = 8'h73 == _t_T_50[15:8] ? 8'h8f : _GEN_6258; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6260 = 8'h74 == _t_T_50[15:8] ? 8'h92 : _GEN_6259; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6261 = 8'h75 == _t_T_50[15:8] ? 8'h9d : _GEN_6260; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6262 = 8'h76 == _t_T_50[15:8] ? 8'h38 : _GEN_6261; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6263 = 8'h77 == _t_T_50[15:8] ? 8'hf5 : _GEN_6262; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6264 = 8'h78 == _t_T_50[15:8] ? 8'hbc : _GEN_6263; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6265 = 8'h79 == _t_T_50[15:8] ? 8'hb6 : _GEN_6264; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6266 = 8'h7a == _t_T_50[15:8] ? 8'hda : _GEN_6265; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6267 = 8'h7b == _t_T_50[15:8] ? 8'h21 : _GEN_6266; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6268 = 8'h7c == _t_T_50[15:8] ? 8'h10 : _GEN_6267; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6269 = 8'h7d == _t_T_50[15:8] ? 8'hff : _GEN_6268; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6270 = 8'h7e == _t_T_50[15:8] ? 8'hf3 : _GEN_6269; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6271 = 8'h7f == _t_T_50[15:8] ? 8'hd2 : _GEN_6270; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6272 = 8'h80 == _t_T_50[15:8] ? 8'hcd : _GEN_6271; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6273 = 8'h81 == _t_T_50[15:8] ? 8'hc : _GEN_6272; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6274 = 8'h82 == _t_T_50[15:8] ? 8'h13 : _GEN_6273; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6275 = 8'h83 == _t_T_50[15:8] ? 8'hec : _GEN_6274; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6276 = 8'h84 == _t_T_50[15:8] ? 8'h5f : _GEN_6275; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6277 = 8'h85 == _t_T_50[15:8] ? 8'h97 : _GEN_6276; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6278 = 8'h86 == _t_T_50[15:8] ? 8'h44 : _GEN_6277; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6279 = 8'h87 == _t_T_50[15:8] ? 8'h17 : _GEN_6278; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6280 = 8'h88 == _t_T_50[15:8] ? 8'hc4 : _GEN_6279; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6281 = 8'h89 == _t_T_50[15:8] ? 8'ha7 : _GEN_6280; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6282 = 8'h8a == _t_T_50[15:8] ? 8'h7e : _GEN_6281; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6283 = 8'h8b == _t_T_50[15:8] ? 8'h3d : _GEN_6282; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6284 = 8'h8c == _t_T_50[15:8] ? 8'h64 : _GEN_6283; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6285 = 8'h8d == _t_T_50[15:8] ? 8'h5d : _GEN_6284; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6286 = 8'h8e == _t_T_50[15:8] ? 8'h19 : _GEN_6285; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6287 = 8'h8f == _t_T_50[15:8] ? 8'h73 : _GEN_6286; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6288 = 8'h90 == _t_T_50[15:8] ? 8'h60 : _GEN_6287; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6289 = 8'h91 == _t_T_50[15:8] ? 8'h81 : _GEN_6288; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6290 = 8'h92 == _t_T_50[15:8] ? 8'h4f : _GEN_6289; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6291 = 8'h93 == _t_T_50[15:8] ? 8'hdc : _GEN_6290; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6292 = 8'h94 == _t_T_50[15:8] ? 8'h22 : _GEN_6291; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6293 = 8'h95 == _t_T_50[15:8] ? 8'h2a : _GEN_6292; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6294 = 8'h96 == _t_T_50[15:8] ? 8'h90 : _GEN_6293; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6295 = 8'h97 == _t_T_50[15:8] ? 8'h88 : _GEN_6294; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6296 = 8'h98 == _t_T_50[15:8] ? 8'h46 : _GEN_6295; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6297 = 8'h99 == _t_T_50[15:8] ? 8'hee : _GEN_6296; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6298 = 8'h9a == _t_T_50[15:8] ? 8'hb8 : _GEN_6297; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6299 = 8'h9b == _t_T_50[15:8] ? 8'h14 : _GEN_6298; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6300 = 8'h9c == _t_T_50[15:8] ? 8'hde : _GEN_6299; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6301 = 8'h9d == _t_T_50[15:8] ? 8'h5e : _GEN_6300; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6302 = 8'h9e == _t_T_50[15:8] ? 8'hb : _GEN_6301; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6303 = 8'h9f == _t_T_50[15:8] ? 8'hdb : _GEN_6302; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6304 = 8'ha0 == _t_T_50[15:8] ? 8'he0 : _GEN_6303; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6305 = 8'ha1 == _t_T_50[15:8] ? 8'h32 : _GEN_6304; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6306 = 8'ha2 == _t_T_50[15:8] ? 8'h3a : _GEN_6305; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6307 = 8'ha3 == _t_T_50[15:8] ? 8'ha : _GEN_6306; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6308 = 8'ha4 == _t_T_50[15:8] ? 8'h49 : _GEN_6307; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6309 = 8'ha5 == _t_T_50[15:8] ? 8'h6 : _GEN_6308; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6310 = 8'ha6 == _t_T_50[15:8] ? 8'h24 : _GEN_6309; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6311 = 8'ha7 == _t_T_50[15:8] ? 8'h5c : _GEN_6310; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6312 = 8'ha8 == _t_T_50[15:8] ? 8'hc2 : _GEN_6311; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6313 = 8'ha9 == _t_T_50[15:8] ? 8'hd3 : _GEN_6312; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6314 = 8'haa == _t_T_50[15:8] ? 8'hac : _GEN_6313; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6315 = 8'hab == _t_T_50[15:8] ? 8'h62 : _GEN_6314; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6316 = 8'hac == _t_T_50[15:8] ? 8'h91 : _GEN_6315; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6317 = 8'had == _t_T_50[15:8] ? 8'h95 : _GEN_6316; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6318 = 8'hae == _t_T_50[15:8] ? 8'he4 : _GEN_6317; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6319 = 8'haf == _t_T_50[15:8] ? 8'h79 : _GEN_6318; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6320 = 8'hb0 == _t_T_50[15:8] ? 8'he7 : _GEN_6319; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6321 = 8'hb1 == _t_T_50[15:8] ? 8'hc8 : _GEN_6320; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6322 = 8'hb2 == _t_T_50[15:8] ? 8'h37 : _GEN_6321; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6323 = 8'hb3 == _t_T_50[15:8] ? 8'h6d : _GEN_6322; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6324 = 8'hb4 == _t_T_50[15:8] ? 8'h8d : _GEN_6323; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6325 = 8'hb5 == _t_T_50[15:8] ? 8'hd5 : _GEN_6324; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6326 = 8'hb6 == _t_T_50[15:8] ? 8'h4e : _GEN_6325; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6327 = 8'hb7 == _t_T_50[15:8] ? 8'ha9 : _GEN_6326; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6328 = 8'hb8 == _t_T_50[15:8] ? 8'h6c : _GEN_6327; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6329 = 8'hb9 == _t_T_50[15:8] ? 8'h56 : _GEN_6328; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6330 = 8'hba == _t_T_50[15:8] ? 8'hf4 : _GEN_6329; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6331 = 8'hbb == _t_T_50[15:8] ? 8'hea : _GEN_6330; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6332 = 8'hbc == _t_T_50[15:8] ? 8'h65 : _GEN_6331; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6333 = 8'hbd == _t_T_50[15:8] ? 8'h7a : _GEN_6332; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6334 = 8'hbe == _t_T_50[15:8] ? 8'hae : _GEN_6333; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6335 = 8'hbf == _t_T_50[15:8] ? 8'h8 : _GEN_6334; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6336 = 8'hc0 == _t_T_50[15:8] ? 8'hba : _GEN_6335; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6337 = 8'hc1 == _t_T_50[15:8] ? 8'h78 : _GEN_6336; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6338 = 8'hc2 == _t_T_50[15:8] ? 8'h25 : _GEN_6337; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6339 = 8'hc3 == _t_T_50[15:8] ? 8'h2e : _GEN_6338; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6340 = 8'hc4 == _t_T_50[15:8] ? 8'h1c : _GEN_6339; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6341 = 8'hc5 == _t_T_50[15:8] ? 8'ha6 : _GEN_6340; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6342 = 8'hc6 == _t_T_50[15:8] ? 8'hb4 : _GEN_6341; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6343 = 8'hc7 == _t_T_50[15:8] ? 8'hc6 : _GEN_6342; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6344 = 8'hc8 == _t_T_50[15:8] ? 8'he8 : _GEN_6343; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6345 = 8'hc9 == _t_T_50[15:8] ? 8'hdd : _GEN_6344; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6346 = 8'hca == _t_T_50[15:8] ? 8'h74 : _GEN_6345; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6347 = 8'hcb == _t_T_50[15:8] ? 8'h1f : _GEN_6346; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6348 = 8'hcc == _t_T_50[15:8] ? 8'h4b : _GEN_6347; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6349 = 8'hcd == _t_T_50[15:8] ? 8'hbd : _GEN_6348; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6350 = 8'hce == _t_T_50[15:8] ? 8'h8b : _GEN_6349; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6351 = 8'hcf == _t_T_50[15:8] ? 8'h8a : _GEN_6350; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6352 = 8'hd0 == _t_T_50[15:8] ? 8'h70 : _GEN_6351; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6353 = 8'hd1 == _t_T_50[15:8] ? 8'h3e : _GEN_6352; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6354 = 8'hd2 == _t_T_50[15:8] ? 8'hb5 : _GEN_6353; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6355 = 8'hd3 == _t_T_50[15:8] ? 8'h66 : _GEN_6354; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6356 = 8'hd4 == _t_T_50[15:8] ? 8'h48 : _GEN_6355; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6357 = 8'hd5 == _t_T_50[15:8] ? 8'h3 : _GEN_6356; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6358 = 8'hd6 == _t_T_50[15:8] ? 8'hf6 : _GEN_6357; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6359 = 8'hd7 == _t_T_50[15:8] ? 8'he : _GEN_6358; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6360 = 8'hd8 == _t_T_50[15:8] ? 8'h61 : _GEN_6359; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6361 = 8'hd9 == _t_T_50[15:8] ? 8'h35 : _GEN_6360; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6362 = 8'hda == _t_T_50[15:8] ? 8'h57 : _GEN_6361; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6363 = 8'hdb == _t_T_50[15:8] ? 8'hb9 : _GEN_6362; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6364 = 8'hdc == _t_T_50[15:8] ? 8'h86 : _GEN_6363; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6365 = 8'hdd == _t_T_50[15:8] ? 8'hc1 : _GEN_6364; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6366 = 8'hde == _t_T_50[15:8] ? 8'h1d : _GEN_6365; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6367 = 8'hdf == _t_T_50[15:8] ? 8'h9e : _GEN_6366; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6368 = 8'he0 == _t_T_50[15:8] ? 8'he1 : _GEN_6367; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6369 = 8'he1 == _t_T_50[15:8] ? 8'hf8 : _GEN_6368; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6370 = 8'he2 == _t_T_50[15:8] ? 8'h98 : _GEN_6369; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6371 = 8'he3 == _t_T_50[15:8] ? 8'h11 : _GEN_6370; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6372 = 8'he4 == _t_T_50[15:8] ? 8'h69 : _GEN_6371; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6373 = 8'he5 == _t_T_50[15:8] ? 8'hd9 : _GEN_6372; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6374 = 8'he6 == _t_T_50[15:8] ? 8'h8e : _GEN_6373; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6375 = 8'he7 == _t_T_50[15:8] ? 8'h94 : _GEN_6374; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6376 = 8'he8 == _t_T_50[15:8] ? 8'h9b : _GEN_6375; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6377 = 8'he9 == _t_T_50[15:8] ? 8'h1e : _GEN_6376; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6378 = 8'hea == _t_T_50[15:8] ? 8'h87 : _GEN_6377; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6379 = 8'heb == _t_T_50[15:8] ? 8'he9 : _GEN_6378; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6380 = 8'hec == _t_T_50[15:8] ? 8'hce : _GEN_6379; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6381 = 8'hed == _t_T_50[15:8] ? 8'h55 : _GEN_6380; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6382 = 8'hee == _t_T_50[15:8] ? 8'h28 : _GEN_6381; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6383 = 8'hef == _t_T_50[15:8] ? 8'hdf : _GEN_6382; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6384 = 8'hf0 == _t_T_50[15:8] ? 8'h8c : _GEN_6383; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6385 = 8'hf1 == _t_T_50[15:8] ? 8'ha1 : _GEN_6384; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6386 = 8'hf2 == _t_T_50[15:8] ? 8'h89 : _GEN_6385; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6387 = 8'hf3 == _t_T_50[15:8] ? 8'hd : _GEN_6386; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6388 = 8'hf4 == _t_T_50[15:8] ? 8'hbf : _GEN_6387; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6389 = 8'hf5 == _t_T_50[15:8] ? 8'he6 : _GEN_6388; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6390 = 8'hf6 == _t_T_50[15:8] ? 8'h42 : _GEN_6389; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6391 = 8'hf7 == _t_T_50[15:8] ? 8'h68 : _GEN_6390; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6392 = 8'hf8 == _t_T_50[15:8] ? 8'h41 : _GEN_6391; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6393 = 8'hf9 == _t_T_50[15:8] ? 8'h99 : _GEN_6392; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6394 = 8'hfa == _t_T_50[15:8] ? 8'h2d : _GEN_6393; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6395 = 8'hfb == _t_T_50[15:8] ? 8'hf : _GEN_6394; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6396 = 8'hfc == _t_T_50[15:8] ? 8'hb0 : _GEN_6395; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6397 = 8'hfd == _t_T_50[15:8] ? 8'h54 : _GEN_6396; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6398 = 8'hfe == _t_T_50[15:8] ? 8'hbb : _GEN_6397; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6399 = 8'hff == _t_T_50[15:8] ? 8'h16 : _GEN_6398; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6401 = 8'h1 == _t_T_50[7:0] ? 8'h7c : 8'h63; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6402 = 8'h2 == _t_T_50[7:0] ? 8'h77 : _GEN_6401; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6403 = 8'h3 == _t_T_50[7:0] ? 8'h7b : _GEN_6402; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6404 = 8'h4 == _t_T_50[7:0] ? 8'hf2 : _GEN_6403; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6405 = 8'h5 == _t_T_50[7:0] ? 8'h6b : _GEN_6404; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6406 = 8'h6 == _t_T_50[7:0] ? 8'h6f : _GEN_6405; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6407 = 8'h7 == _t_T_50[7:0] ? 8'hc5 : _GEN_6406; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6408 = 8'h8 == _t_T_50[7:0] ? 8'h30 : _GEN_6407; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6409 = 8'h9 == _t_T_50[7:0] ? 8'h1 : _GEN_6408; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6410 = 8'ha == _t_T_50[7:0] ? 8'h67 : _GEN_6409; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6411 = 8'hb == _t_T_50[7:0] ? 8'h2b : _GEN_6410; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6412 = 8'hc == _t_T_50[7:0] ? 8'hfe : _GEN_6411; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6413 = 8'hd == _t_T_50[7:0] ? 8'hd7 : _GEN_6412; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6414 = 8'he == _t_T_50[7:0] ? 8'hab : _GEN_6413; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6415 = 8'hf == _t_T_50[7:0] ? 8'h76 : _GEN_6414; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6416 = 8'h10 == _t_T_50[7:0] ? 8'hca : _GEN_6415; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6417 = 8'h11 == _t_T_50[7:0] ? 8'h82 : _GEN_6416; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6418 = 8'h12 == _t_T_50[7:0] ? 8'hc9 : _GEN_6417; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6419 = 8'h13 == _t_T_50[7:0] ? 8'h7d : _GEN_6418; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6420 = 8'h14 == _t_T_50[7:0] ? 8'hfa : _GEN_6419; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6421 = 8'h15 == _t_T_50[7:0] ? 8'h59 : _GEN_6420; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6422 = 8'h16 == _t_T_50[7:0] ? 8'h47 : _GEN_6421; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6423 = 8'h17 == _t_T_50[7:0] ? 8'hf0 : _GEN_6422; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6424 = 8'h18 == _t_T_50[7:0] ? 8'had : _GEN_6423; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6425 = 8'h19 == _t_T_50[7:0] ? 8'hd4 : _GEN_6424; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6426 = 8'h1a == _t_T_50[7:0] ? 8'ha2 : _GEN_6425; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6427 = 8'h1b == _t_T_50[7:0] ? 8'haf : _GEN_6426; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6428 = 8'h1c == _t_T_50[7:0] ? 8'h9c : _GEN_6427; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6429 = 8'h1d == _t_T_50[7:0] ? 8'ha4 : _GEN_6428; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6430 = 8'h1e == _t_T_50[7:0] ? 8'h72 : _GEN_6429; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6431 = 8'h1f == _t_T_50[7:0] ? 8'hc0 : _GEN_6430; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6432 = 8'h20 == _t_T_50[7:0] ? 8'hb7 : _GEN_6431; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6433 = 8'h21 == _t_T_50[7:0] ? 8'hfd : _GEN_6432; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6434 = 8'h22 == _t_T_50[7:0] ? 8'h93 : _GEN_6433; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6435 = 8'h23 == _t_T_50[7:0] ? 8'h26 : _GEN_6434; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6436 = 8'h24 == _t_T_50[7:0] ? 8'h36 : _GEN_6435; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6437 = 8'h25 == _t_T_50[7:0] ? 8'h3f : _GEN_6436; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6438 = 8'h26 == _t_T_50[7:0] ? 8'hf7 : _GEN_6437; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6439 = 8'h27 == _t_T_50[7:0] ? 8'hcc : _GEN_6438; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6440 = 8'h28 == _t_T_50[7:0] ? 8'h34 : _GEN_6439; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6441 = 8'h29 == _t_T_50[7:0] ? 8'ha5 : _GEN_6440; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6442 = 8'h2a == _t_T_50[7:0] ? 8'he5 : _GEN_6441; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6443 = 8'h2b == _t_T_50[7:0] ? 8'hf1 : _GEN_6442; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6444 = 8'h2c == _t_T_50[7:0] ? 8'h71 : _GEN_6443; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6445 = 8'h2d == _t_T_50[7:0] ? 8'hd8 : _GEN_6444; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6446 = 8'h2e == _t_T_50[7:0] ? 8'h31 : _GEN_6445; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6447 = 8'h2f == _t_T_50[7:0] ? 8'h15 : _GEN_6446; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6448 = 8'h30 == _t_T_50[7:0] ? 8'h4 : _GEN_6447; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6449 = 8'h31 == _t_T_50[7:0] ? 8'hc7 : _GEN_6448; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6450 = 8'h32 == _t_T_50[7:0] ? 8'h23 : _GEN_6449; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6451 = 8'h33 == _t_T_50[7:0] ? 8'hc3 : _GEN_6450; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6452 = 8'h34 == _t_T_50[7:0] ? 8'h18 : _GEN_6451; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6453 = 8'h35 == _t_T_50[7:0] ? 8'h96 : _GEN_6452; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6454 = 8'h36 == _t_T_50[7:0] ? 8'h5 : _GEN_6453; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6455 = 8'h37 == _t_T_50[7:0] ? 8'h9a : _GEN_6454; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6456 = 8'h38 == _t_T_50[7:0] ? 8'h7 : _GEN_6455; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6457 = 8'h39 == _t_T_50[7:0] ? 8'h12 : _GEN_6456; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6458 = 8'h3a == _t_T_50[7:0] ? 8'h80 : _GEN_6457; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6459 = 8'h3b == _t_T_50[7:0] ? 8'he2 : _GEN_6458; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6460 = 8'h3c == _t_T_50[7:0] ? 8'heb : _GEN_6459; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6461 = 8'h3d == _t_T_50[7:0] ? 8'h27 : _GEN_6460; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6462 = 8'h3e == _t_T_50[7:0] ? 8'hb2 : _GEN_6461; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6463 = 8'h3f == _t_T_50[7:0] ? 8'h75 : _GEN_6462; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6464 = 8'h40 == _t_T_50[7:0] ? 8'h9 : _GEN_6463; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6465 = 8'h41 == _t_T_50[7:0] ? 8'h83 : _GEN_6464; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6466 = 8'h42 == _t_T_50[7:0] ? 8'h2c : _GEN_6465; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6467 = 8'h43 == _t_T_50[7:0] ? 8'h1a : _GEN_6466; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6468 = 8'h44 == _t_T_50[7:0] ? 8'h1b : _GEN_6467; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6469 = 8'h45 == _t_T_50[7:0] ? 8'h6e : _GEN_6468; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6470 = 8'h46 == _t_T_50[7:0] ? 8'h5a : _GEN_6469; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6471 = 8'h47 == _t_T_50[7:0] ? 8'ha0 : _GEN_6470; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6472 = 8'h48 == _t_T_50[7:0] ? 8'h52 : _GEN_6471; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6473 = 8'h49 == _t_T_50[7:0] ? 8'h3b : _GEN_6472; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6474 = 8'h4a == _t_T_50[7:0] ? 8'hd6 : _GEN_6473; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6475 = 8'h4b == _t_T_50[7:0] ? 8'hb3 : _GEN_6474; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6476 = 8'h4c == _t_T_50[7:0] ? 8'h29 : _GEN_6475; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6477 = 8'h4d == _t_T_50[7:0] ? 8'he3 : _GEN_6476; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6478 = 8'h4e == _t_T_50[7:0] ? 8'h2f : _GEN_6477; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6479 = 8'h4f == _t_T_50[7:0] ? 8'h84 : _GEN_6478; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6480 = 8'h50 == _t_T_50[7:0] ? 8'h53 : _GEN_6479; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6481 = 8'h51 == _t_T_50[7:0] ? 8'hd1 : _GEN_6480; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6482 = 8'h52 == _t_T_50[7:0] ? 8'h0 : _GEN_6481; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6483 = 8'h53 == _t_T_50[7:0] ? 8'hed : _GEN_6482; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6484 = 8'h54 == _t_T_50[7:0] ? 8'h20 : _GEN_6483; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6485 = 8'h55 == _t_T_50[7:0] ? 8'hfc : _GEN_6484; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6486 = 8'h56 == _t_T_50[7:0] ? 8'hb1 : _GEN_6485; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6487 = 8'h57 == _t_T_50[7:0] ? 8'h5b : _GEN_6486; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6488 = 8'h58 == _t_T_50[7:0] ? 8'h6a : _GEN_6487; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6489 = 8'h59 == _t_T_50[7:0] ? 8'hcb : _GEN_6488; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6490 = 8'h5a == _t_T_50[7:0] ? 8'hbe : _GEN_6489; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6491 = 8'h5b == _t_T_50[7:0] ? 8'h39 : _GEN_6490; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6492 = 8'h5c == _t_T_50[7:0] ? 8'h4a : _GEN_6491; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6493 = 8'h5d == _t_T_50[7:0] ? 8'h4c : _GEN_6492; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6494 = 8'h5e == _t_T_50[7:0] ? 8'h58 : _GEN_6493; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6495 = 8'h5f == _t_T_50[7:0] ? 8'hcf : _GEN_6494; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6496 = 8'h60 == _t_T_50[7:0] ? 8'hd0 : _GEN_6495; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6497 = 8'h61 == _t_T_50[7:0] ? 8'hef : _GEN_6496; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6498 = 8'h62 == _t_T_50[7:0] ? 8'haa : _GEN_6497; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6499 = 8'h63 == _t_T_50[7:0] ? 8'hfb : _GEN_6498; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6500 = 8'h64 == _t_T_50[7:0] ? 8'h43 : _GEN_6499; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6501 = 8'h65 == _t_T_50[7:0] ? 8'h4d : _GEN_6500; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6502 = 8'h66 == _t_T_50[7:0] ? 8'h33 : _GEN_6501; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6503 = 8'h67 == _t_T_50[7:0] ? 8'h85 : _GEN_6502; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6504 = 8'h68 == _t_T_50[7:0] ? 8'h45 : _GEN_6503; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6505 = 8'h69 == _t_T_50[7:0] ? 8'hf9 : _GEN_6504; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6506 = 8'h6a == _t_T_50[7:0] ? 8'h2 : _GEN_6505; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6507 = 8'h6b == _t_T_50[7:0] ? 8'h7f : _GEN_6506; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6508 = 8'h6c == _t_T_50[7:0] ? 8'h50 : _GEN_6507; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6509 = 8'h6d == _t_T_50[7:0] ? 8'h3c : _GEN_6508; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6510 = 8'h6e == _t_T_50[7:0] ? 8'h9f : _GEN_6509; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6511 = 8'h6f == _t_T_50[7:0] ? 8'ha8 : _GEN_6510; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6512 = 8'h70 == _t_T_50[7:0] ? 8'h51 : _GEN_6511; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6513 = 8'h71 == _t_T_50[7:0] ? 8'ha3 : _GEN_6512; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6514 = 8'h72 == _t_T_50[7:0] ? 8'h40 : _GEN_6513; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6515 = 8'h73 == _t_T_50[7:0] ? 8'h8f : _GEN_6514; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6516 = 8'h74 == _t_T_50[7:0] ? 8'h92 : _GEN_6515; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6517 = 8'h75 == _t_T_50[7:0] ? 8'h9d : _GEN_6516; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6518 = 8'h76 == _t_T_50[7:0] ? 8'h38 : _GEN_6517; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6519 = 8'h77 == _t_T_50[7:0] ? 8'hf5 : _GEN_6518; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6520 = 8'h78 == _t_T_50[7:0] ? 8'hbc : _GEN_6519; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6521 = 8'h79 == _t_T_50[7:0] ? 8'hb6 : _GEN_6520; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6522 = 8'h7a == _t_T_50[7:0] ? 8'hda : _GEN_6521; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6523 = 8'h7b == _t_T_50[7:0] ? 8'h21 : _GEN_6522; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6524 = 8'h7c == _t_T_50[7:0] ? 8'h10 : _GEN_6523; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6525 = 8'h7d == _t_T_50[7:0] ? 8'hff : _GEN_6524; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6526 = 8'h7e == _t_T_50[7:0] ? 8'hf3 : _GEN_6525; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6527 = 8'h7f == _t_T_50[7:0] ? 8'hd2 : _GEN_6526; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6528 = 8'h80 == _t_T_50[7:0] ? 8'hcd : _GEN_6527; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6529 = 8'h81 == _t_T_50[7:0] ? 8'hc : _GEN_6528; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6530 = 8'h82 == _t_T_50[7:0] ? 8'h13 : _GEN_6529; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6531 = 8'h83 == _t_T_50[7:0] ? 8'hec : _GEN_6530; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6532 = 8'h84 == _t_T_50[7:0] ? 8'h5f : _GEN_6531; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6533 = 8'h85 == _t_T_50[7:0] ? 8'h97 : _GEN_6532; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6534 = 8'h86 == _t_T_50[7:0] ? 8'h44 : _GEN_6533; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6535 = 8'h87 == _t_T_50[7:0] ? 8'h17 : _GEN_6534; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6536 = 8'h88 == _t_T_50[7:0] ? 8'hc4 : _GEN_6535; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6537 = 8'h89 == _t_T_50[7:0] ? 8'ha7 : _GEN_6536; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6538 = 8'h8a == _t_T_50[7:0] ? 8'h7e : _GEN_6537; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6539 = 8'h8b == _t_T_50[7:0] ? 8'h3d : _GEN_6538; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6540 = 8'h8c == _t_T_50[7:0] ? 8'h64 : _GEN_6539; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6541 = 8'h8d == _t_T_50[7:0] ? 8'h5d : _GEN_6540; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6542 = 8'h8e == _t_T_50[7:0] ? 8'h19 : _GEN_6541; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6543 = 8'h8f == _t_T_50[7:0] ? 8'h73 : _GEN_6542; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6544 = 8'h90 == _t_T_50[7:0] ? 8'h60 : _GEN_6543; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6545 = 8'h91 == _t_T_50[7:0] ? 8'h81 : _GEN_6544; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6546 = 8'h92 == _t_T_50[7:0] ? 8'h4f : _GEN_6545; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6547 = 8'h93 == _t_T_50[7:0] ? 8'hdc : _GEN_6546; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6548 = 8'h94 == _t_T_50[7:0] ? 8'h22 : _GEN_6547; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6549 = 8'h95 == _t_T_50[7:0] ? 8'h2a : _GEN_6548; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6550 = 8'h96 == _t_T_50[7:0] ? 8'h90 : _GEN_6549; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6551 = 8'h97 == _t_T_50[7:0] ? 8'h88 : _GEN_6550; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6552 = 8'h98 == _t_T_50[7:0] ? 8'h46 : _GEN_6551; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6553 = 8'h99 == _t_T_50[7:0] ? 8'hee : _GEN_6552; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6554 = 8'h9a == _t_T_50[7:0] ? 8'hb8 : _GEN_6553; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6555 = 8'h9b == _t_T_50[7:0] ? 8'h14 : _GEN_6554; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6556 = 8'h9c == _t_T_50[7:0] ? 8'hde : _GEN_6555; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6557 = 8'h9d == _t_T_50[7:0] ? 8'h5e : _GEN_6556; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6558 = 8'h9e == _t_T_50[7:0] ? 8'hb : _GEN_6557; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6559 = 8'h9f == _t_T_50[7:0] ? 8'hdb : _GEN_6558; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6560 = 8'ha0 == _t_T_50[7:0] ? 8'he0 : _GEN_6559; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6561 = 8'ha1 == _t_T_50[7:0] ? 8'h32 : _GEN_6560; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6562 = 8'ha2 == _t_T_50[7:0] ? 8'h3a : _GEN_6561; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6563 = 8'ha3 == _t_T_50[7:0] ? 8'ha : _GEN_6562; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6564 = 8'ha4 == _t_T_50[7:0] ? 8'h49 : _GEN_6563; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6565 = 8'ha5 == _t_T_50[7:0] ? 8'h6 : _GEN_6564; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6566 = 8'ha6 == _t_T_50[7:0] ? 8'h24 : _GEN_6565; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6567 = 8'ha7 == _t_T_50[7:0] ? 8'h5c : _GEN_6566; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6568 = 8'ha8 == _t_T_50[7:0] ? 8'hc2 : _GEN_6567; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6569 = 8'ha9 == _t_T_50[7:0] ? 8'hd3 : _GEN_6568; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6570 = 8'haa == _t_T_50[7:0] ? 8'hac : _GEN_6569; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6571 = 8'hab == _t_T_50[7:0] ? 8'h62 : _GEN_6570; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6572 = 8'hac == _t_T_50[7:0] ? 8'h91 : _GEN_6571; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6573 = 8'had == _t_T_50[7:0] ? 8'h95 : _GEN_6572; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6574 = 8'hae == _t_T_50[7:0] ? 8'he4 : _GEN_6573; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6575 = 8'haf == _t_T_50[7:0] ? 8'h79 : _GEN_6574; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6576 = 8'hb0 == _t_T_50[7:0] ? 8'he7 : _GEN_6575; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6577 = 8'hb1 == _t_T_50[7:0] ? 8'hc8 : _GEN_6576; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6578 = 8'hb2 == _t_T_50[7:0] ? 8'h37 : _GEN_6577; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6579 = 8'hb3 == _t_T_50[7:0] ? 8'h6d : _GEN_6578; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6580 = 8'hb4 == _t_T_50[7:0] ? 8'h8d : _GEN_6579; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6581 = 8'hb5 == _t_T_50[7:0] ? 8'hd5 : _GEN_6580; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6582 = 8'hb6 == _t_T_50[7:0] ? 8'h4e : _GEN_6581; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6583 = 8'hb7 == _t_T_50[7:0] ? 8'ha9 : _GEN_6582; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6584 = 8'hb8 == _t_T_50[7:0] ? 8'h6c : _GEN_6583; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6585 = 8'hb9 == _t_T_50[7:0] ? 8'h56 : _GEN_6584; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6586 = 8'hba == _t_T_50[7:0] ? 8'hf4 : _GEN_6585; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6587 = 8'hbb == _t_T_50[7:0] ? 8'hea : _GEN_6586; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6588 = 8'hbc == _t_T_50[7:0] ? 8'h65 : _GEN_6587; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6589 = 8'hbd == _t_T_50[7:0] ? 8'h7a : _GEN_6588; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6590 = 8'hbe == _t_T_50[7:0] ? 8'hae : _GEN_6589; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6591 = 8'hbf == _t_T_50[7:0] ? 8'h8 : _GEN_6590; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6592 = 8'hc0 == _t_T_50[7:0] ? 8'hba : _GEN_6591; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6593 = 8'hc1 == _t_T_50[7:0] ? 8'h78 : _GEN_6592; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6594 = 8'hc2 == _t_T_50[7:0] ? 8'h25 : _GEN_6593; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6595 = 8'hc3 == _t_T_50[7:0] ? 8'h2e : _GEN_6594; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6596 = 8'hc4 == _t_T_50[7:0] ? 8'h1c : _GEN_6595; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6597 = 8'hc5 == _t_T_50[7:0] ? 8'ha6 : _GEN_6596; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6598 = 8'hc6 == _t_T_50[7:0] ? 8'hb4 : _GEN_6597; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6599 = 8'hc7 == _t_T_50[7:0] ? 8'hc6 : _GEN_6598; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6600 = 8'hc8 == _t_T_50[7:0] ? 8'he8 : _GEN_6599; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6601 = 8'hc9 == _t_T_50[7:0] ? 8'hdd : _GEN_6600; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6602 = 8'hca == _t_T_50[7:0] ? 8'h74 : _GEN_6601; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6603 = 8'hcb == _t_T_50[7:0] ? 8'h1f : _GEN_6602; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6604 = 8'hcc == _t_T_50[7:0] ? 8'h4b : _GEN_6603; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6605 = 8'hcd == _t_T_50[7:0] ? 8'hbd : _GEN_6604; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6606 = 8'hce == _t_T_50[7:0] ? 8'h8b : _GEN_6605; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6607 = 8'hcf == _t_T_50[7:0] ? 8'h8a : _GEN_6606; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6608 = 8'hd0 == _t_T_50[7:0] ? 8'h70 : _GEN_6607; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6609 = 8'hd1 == _t_T_50[7:0] ? 8'h3e : _GEN_6608; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6610 = 8'hd2 == _t_T_50[7:0] ? 8'hb5 : _GEN_6609; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6611 = 8'hd3 == _t_T_50[7:0] ? 8'h66 : _GEN_6610; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6612 = 8'hd4 == _t_T_50[7:0] ? 8'h48 : _GEN_6611; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6613 = 8'hd5 == _t_T_50[7:0] ? 8'h3 : _GEN_6612; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6614 = 8'hd6 == _t_T_50[7:0] ? 8'hf6 : _GEN_6613; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6615 = 8'hd7 == _t_T_50[7:0] ? 8'he : _GEN_6614; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6616 = 8'hd8 == _t_T_50[7:0] ? 8'h61 : _GEN_6615; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6617 = 8'hd9 == _t_T_50[7:0] ? 8'h35 : _GEN_6616; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6618 = 8'hda == _t_T_50[7:0] ? 8'h57 : _GEN_6617; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6619 = 8'hdb == _t_T_50[7:0] ? 8'hb9 : _GEN_6618; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6620 = 8'hdc == _t_T_50[7:0] ? 8'h86 : _GEN_6619; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6621 = 8'hdd == _t_T_50[7:0] ? 8'hc1 : _GEN_6620; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6622 = 8'hde == _t_T_50[7:0] ? 8'h1d : _GEN_6621; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6623 = 8'hdf == _t_T_50[7:0] ? 8'h9e : _GEN_6622; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6624 = 8'he0 == _t_T_50[7:0] ? 8'he1 : _GEN_6623; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6625 = 8'he1 == _t_T_50[7:0] ? 8'hf8 : _GEN_6624; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6626 = 8'he2 == _t_T_50[7:0] ? 8'h98 : _GEN_6625; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6627 = 8'he3 == _t_T_50[7:0] ? 8'h11 : _GEN_6626; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6628 = 8'he4 == _t_T_50[7:0] ? 8'h69 : _GEN_6627; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6629 = 8'he5 == _t_T_50[7:0] ? 8'hd9 : _GEN_6628; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6630 = 8'he6 == _t_T_50[7:0] ? 8'h8e : _GEN_6629; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6631 = 8'he7 == _t_T_50[7:0] ? 8'h94 : _GEN_6630; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6632 = 8'he8 == _t_T_50[7:0] ? 8'h9b : _GEN_6631; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6633 = 8'he9 == _t_T_50[7:0] ? 8'h1e : _GEN_6632; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6634 = 8'hea == _t_T_50[7:0] ? 8'h87 : _GEN_6633; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6635 = 8'heb == _t_T_50[7:0] ? 8'he9 : _GEN_6634; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6636 = 8'hec == _t_T_50[7:0] ? 8'hce : _GEN_6635; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6637 = 8'hed == _t_T_50[7:0] ? 8'h55 : _GEN_6636; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6638 = 8'hee == _t_T_50[7:0] ? 8'h28 : _GEN_6637; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6639 = 8'hef == _t_T_50[7:0] ? 8'hdf : _GEN_6638; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6640 = 8'hf0 == _t_T_50[7:0] ? 8'h8c : _GEN_6639; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6641 = 8'hf1 == _t_T_50[7:0] ? 8'ha1 : _GEN_6640; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6642 = 8'hf2 == _t_T_50[7:0] ? 8'h89 : _GEN_6641; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6643 = 8'hf3 == _t_T_50[7:0] ? 8'hd : _GEN_6642; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6644 = 8'hf4 == _t_T_50[7:0] ? 8'hbf : _GEN_6643; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6645 = 8'hf5 == _t_T_50[7:0] ? 8'he6 : _GEN_6644; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6646 = 8'hf6 == _t_T_50[7:0] ? 8'h42 : _GEN_6645; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6647 = 8'hf7 == _t_T_50[7:0] ? 8'h68 : _GEN_6646; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6648 = 8'hf8 == _t_T_50[7:0] ? 8'h41 : _GEN_6647; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6649 = 8'hf9 == _t_T_50[7:0] ? 8'h99 : _GEN_6648; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6650 = 8'hfa == _t_T_50[7:0] ? 8'h2d : _GEN_6649; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6651 = 8'hfb == _t_T_50[7:0] ? 8'hf : _GEN_6650; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6652 = 8'hfc == _t_T_50[7:0] ? 8'hb0 : _GEN_6651; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6653 = 8'hfd == _t_T_50[7:0] ? 8'h54 : _GEN_6652; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6654 = 8'hfe == _t_T_50[7:0] ? 8'hbb : _GEN_6653; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6655 = 8'hff == _t_T_50[7:0] ? 8'h16 : _GEN_6654; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6657 = 8'h1 == _t_T_50[31:24] ? 8'h7c : 8'h63; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6658 = 8'h2 == _t_T_50[31:24] ? 8'h77 : _GEN_6657; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6659 = 8'h3 == _t_T_50[31:24] ? 8'h7b : _GEN_6658; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6660 = 8'h4 == _t_T_50[31:24] ? 8'hf2 : _GEN_6659; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6661 = 8'h5 == _t_T_50[31:24] ? 8'h6b : _GEN_6660; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6662 = 8'h6 == _t_T_50[31:24] ? 8'h6f : _GEN_6661; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6663 = 8'h7 == _t_T_50[31:24] ? 8'hc5 : _GEN_6662; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6664 = 8'h8 == _t_T_50[31:24] ? 8'h30 : _GEN_6663; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6665 = 8'h9 == _t_T_50[31:24] ? 8'h1 : _GEN_6664; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6666 = 8'ha == _t_T_50[31:24] ? 8'h67 : _GEN_6665; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6667 = 8'hb == _t_T_50[31:24] ? 8'h2b : _GEN_6666; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6668 = 8'hc == _t_T_50[31:24] ? 8'hfe : _GEN_6667; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6669 = 8'hd == _t_T_50[31:24] ? 8'hd7 : _GEN_6668; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6670 = 8'he == _t_T_50[31:24] ? 8'hab : _GEN_6669; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6671 = 8'hf == _t_T_50[31:24] ? 8'h76 : _GEN_6670; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6672 = 8'h10 == _t_T_50[31:24] ? 8'hca : _GEN_6671; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6673 = 8'h11 == _t_T_50[31:24] ? 8'h82 : _GEN_6672; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6674 = 8'h12 == _t_T_50[31:24] ? 8'hc9 : _GEN_6673; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6675 = 8'h13 == _t_T_50[31:24] ? 8'h7d : _GEN_6674; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6676 = 8'h14 == _t_T_50[31:24] ? 8'hfa : _GEN_6675; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6677 = 8'h15 == _t_T_50[31:24] ? 8'h59 : _GEN_6676; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6678 = 8'h16 == _t_T_50[31:24] ? 8'h47 : _GEN_6677; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6679 = 8'h17 == _t_T_50[31:24] ? 8'hf0 : _GEN_6678; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6680 = 8'h18 == _t_T_50[31:24] ? 8'had : _GEN_6679; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6681 = 8'h19 == _t_T_50[31:24] ? 8'hd4 : _GEN_6680; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6682 = 8'h1a == _t_T_50[31:24] ? 8'ha2 : _GEN_6681; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6683 = 8'h1b == _t_T_50[31:24] ? 8'haf : _GEN_6682; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6684 = 8'h1c == _t_T_50[31:24] ? 8'h9c : _GEN_6683; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6685 = 8'h1d == _t_T_50[31:24] ? 8'ha4 : _GEN_6684; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6686 = 8'h1e == _t_T_50[31:24] ? 8'h72 : _GEN_6685; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6687 = 8'h1f == _t_T_50[31:24] ? 8'hc0 : _GEN_6686; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6688 = 8'h20 == _t_T_50[31:24] ? 8'hb7 : _GEN_6687; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6689 = 8'h21 == _t_T_50[31:24] ? 8'hfd : _GEN_6688; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6690 = 8'h22 == _t_T_50[31:24] ? 8'h93 : _GEN_6689; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6691 = 8'h23 == _t_T_50[31:24] ? 8'h26 : _GEN_6690; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6692 = 8'h24 == _t_T_50[31:24] ? 8'h36 : _GEN_6691; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6693 = 8'h25 == _t_T_50[31:24] ? 8'h3f : _GEN_6692; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6694 = 8'h26 == _t_T_50[31:24] ? 8'hf7 : _GEN_6693; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6695 = 8'h27 == _t_T_50[31:24] ? 8'hcc : _GEN_6694; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6696 = 8'h28 == _t_T_50[31:24] ? 8'h34 : _GEN_6695; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6697 = 8'h29 == _t_T_50[31:24] ? 8'ha5 : _GEN_6696; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6698 = 8'h2a == _t_T_50[31:24] ? 8'he5 : _GEN_6697; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6699 = 8'h2b == _t_T_50[31:24] ? 8'hf1 : _GEN_6698; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6700 = 8'h2c == _t_T_50[31:24] ? 8'h71 : _GEN_6699; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6701 = 8'h2d == _t_T_50[31:24] ? 8'hd8 : _GEN_6700; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6702 = 8'h2e == _t_T_50[31:24] ? 8'h31 : _GEN_6701; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6703 = 8'h2f == _t_T_50[31:24] ? 8'h15 : _GEN_6702; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6704 = 8'h30 == _t_T_50[31:24] ? 8'h4 : _GEN_6703; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6705 = 8'h31 == _t_T_50[31:24] ? 8'hc7 : _GEN_6704; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6706 = 8'h32 == _t_T_50[31:24] ? 8'h23 : _GEN_6705; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6707 = 8'h33 == _t_T_50[31:24] ? 8'hc3 : _GEN_6706; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6708 = 8'h34 == _t_T_50[31:24] ? 8'h18 : _GEN_6707; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6709 = 8'h35 == _t_T_50[31:24] ? 8'h96 : _GEN_6708; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6710 = 8'h36 == _t_T_50[31:24] ? 8'h5 : _GEN_6709; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6711 = 8'h37 == _t_T_50[31:24] ? 8'h9a : _GEN_6710; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6712 = 8'h38 == _t_T_50[31:24] ? 8'h7 : _GEN_6711; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6713 = 8'h39 == _t_T_50[31:24] ? 8'h12 : _GEN_6712; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6714 = 8'h3a == _t_T_50[31:24] ? 8'h80 : _GEN_6713; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6715 = 8'h3b == _t_T_50[31:24] ? 8'he2 : _GEN_6714; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6716 = 8'h3c == _t_T_50[31:24] ? 8'heb : _GEN_6715; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6717 = 8'h3d == _t_T_50[31:24] ? 8'h27 : _GEN_6716; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6718 = 8'h3e == _t_T_50[31:24] ? 8'hb2 : _GEN_6717; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6719 = 8'h3f == _t_T_50[31:24] ? 8'h75 : _GEN_6718; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6720 = 8'h40 == _t_T_50[31:24] ? 8'h9 : _GEN_6719; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6721 = 8'h41 == _t_T_50[31:24] ? 8'h83 : _GEN_6720; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6722 = 8'h42 == _t_T_50[31:24] ? 8'h2c : _GEN_6721; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6723 = 8'h43 == _t_T_50[31:24] ? 8'h1a : _GEN_6722; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6724 = 8'h44 == _t_T_50[31:24] ? 8'h1b : _GEN_6723; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6725 = 8'h45 == _t_T_50[31:24] ? 8'h6e : _GEN_6724; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6726 = 8'h46 == _t_T_50[31:24] ? 8'h5a : _GEN_6725; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6727 = 8'h47 == _t_T_50[31:24] ? 8'ha0 : _GEN_6726; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6728 = 8'h48 == _t_T_50[31:24] ? 8'h52 : _GEN_6727; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6729 = 8'h49 == _t_T_50[31:24] ? 8'h3b : _GEN_6728; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6730 = 8'h4a == _t_T_50[31:24] ? 8'hd6 : _GEN_6729; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6731 = 8'h4b == _t_T_50[31:24] ? 8'hb3 : _GEN_6730; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6732 = 8'h4c == _t_T_50[31:24] ? 8'h29 : _GEN_6731; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6733 = 8'h4d == _t_T_50[31:24] ? 8'he3 : _GEN_6732; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6734 = 8'h4e == _t_T_50[31:24] ? 8'h2f : _GEN_6733; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6735 = 8'h4f == _t_T_50[31:24] ? 8'h84 : _GEN_6734; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6736 = 8'h50 == _t_T_50[31:24] ? 8'h53 : _GEN_6735; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6737 = 8'h51 == _t_T_50[31:24] ? 8'hd1 : _GEN_6736; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6738 = 8'h52 == _t_T_50[31:24] ? 8'h0 : _GEN_6737; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6739 = 8'h53 == _t_T_50[31:24] ? 8'hed : _GEN_6738; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6740 = 8'h54 == _t_T_50[31:24] ? 8'h20 : _GEN_6739; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6741 = 8'h55 == _t_T_50[31:24] ? 8'hfc : _GEN_6740; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6742 = 8'h56 == _t_T_50[31:24] ? 8'hb1 : _GEN_6741; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6743 = 8'h57 == _t_T_50[31:24] ? 8'h5b : _GEN_6742; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6744 = 8'h58 == _t_T_50[31:24] ? 8'h6a : _GEN_6743; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6745 = 8'h59 == _t_T_50[31:24] ? 8'hcb : _GEN_6744; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6746 = 8'h5a == _t_T_50[31:24] ? 8'hbe : _GEN_6745; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6747 = 8'h5b == _t_T_50[31:24] ? 8'h39 : _GEN_6746; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6748 = 8'h5c == _t_T_50[31:24] ? 8'h4a : _GEN_6747; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6749 = 8'h5d == _t_T_50[31:24] ? 8'h4c : _GEN_6748; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6750 = 8'h5e == _t_T_50[31:24] ? 8'h58 : _GEN_6749; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6751 = 8'h5f == _t_T_50[31:24] ? 8'hcf : _GEN_6750; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6752 = 8'h60 == _t_T_50[31:24] ? 8'hd0 : _GEN_6751; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6753 = 8'h61 == _t_T_50[31:24] ? 8'hef : _GEN_6752; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6754 = 8'h62 == _t_T_50[31:24] ? 8'haa : _GEN_6753; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6755 = 8'h63 == _t_T_50[31:24] ? 8'hfb : _GEN_6754; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6756 = 8'h64 == _t_T_50[31:24] ? 8'h43 : _GEN_6755; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6757 = 8'h65 == _t_T_50[31:24] ? 8'h4d : _GEN_6756; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6758 = 8'h66 == _t_T_50[31:24] ? 8'h33 : _GEN_6757; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6759 = 8'h67 == _t_T_50[31:24] ? 8'h85 : _GEN_6758; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6760 = 8'h68 == _t_T_50[31:24] ? 8'h45 : _GEN_6759; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6761 = 8'h69 == _t_T_50[31:24] ? 8'hf9 : _GEN_6760; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6762 = 8'h6a == _t_T_50[31:24] ? 8'h2 : _GEN_6761; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6763 = 8'h6b == _t_T_50[31:24] ? 8'h7f : _GEN_6762; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6764 = 8'h6c == _t_T_50[31:24] ? 8'h50 : _GEN_6763; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6765 = 8'h6d == _t_T_50[31:24] ? 8'h3c : _GEN_6764; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6766 = 8'h6e == _t_T_50[31:24] ? 8'h9f : _GEN_6765; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6767 = 8'h6f == _t_T_50[31:24] ? 8'ha8 : _GEN_6766; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6768 = 8'h70 == _t_T_50[31:24] ? 8'h51 : _GEN_6767; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6769 = 8'h71 == _t_T_50[31:24] ? 8'ha3 : _GEN_6768; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6770 = 8'h72 == _t_T_50[31:24] ? 8'h40 : _GEN_6769; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6771 = 8'h73 == _t_T_50[31:24] ? 8'h8f : _GEN_6770; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6772 = 8'h74 == _t_T_50[31:24] ? 8'h92 : _GEN_6771; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6773 = 8'h75 == _t_T_50[31:24] ? 8'h9d : _GEN_6772; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6774 = 8'h76 == _t_T_50[31:24] ? 8'h38 : _GEN_6773; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6775 = 8'h77 == _t_T_50[31:24] ? 8'hf5 : _GEN_6774; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6776 = 8'h78 == _t_T_50[31:24] ? 8'hbc : _GEN_6775; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6777 = 8'h79 == _t_T_50[31:24] ? 8'hb6 : _GEN_6776; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6778 = 8'h7a == _t_T_50[31:24] ? 8'hda : _GEN_6777; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6779 = 8'h7b == _t_T_50[31:24] ? 8'h21 : _GEN_6778; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6780 = 8'h7c == _t_T_50[31:24] ? 8'h10 : _GEN_6779; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6781 = 8'h7d == _t_T_50[31:24] ? 8'hff : _GEN_6780; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6782 = 8'h7e == _t_T_50[31:24] ? 8'hf3 : _GEN_6781; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6783 = 8'h7f == _t_T_50[31:24] ? 8'hd2 : _GEN_6782; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6784 = 8'h80 == _t_T_50[31:24] ? 8'hcd : _GEN_6783; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6785 = 8'h81 == _t_T_50[31:24] ? 8'hc : _GEN_6784; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6786 = 8'h82 == _t_T_50[31:24] ? 8'h13 : _GEN_6785; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6787 = 8'h83 == _t_T_50[31:24] ? 8'hec : _GEN_6786; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6788 = 8'h84 == _t_T_50[31:24] ? 8'h5f : _GEN_6787; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6789 = 8'h85 == _t_T_50[31:24] ? 8'h97 : _GEN_6788; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6790 = 8'h86 == _t_T_50[31:24] ? 8'h44 : _GEN_6789; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6791 = 8'h87 == _t_T_50[31:24] ? 8'h17 : _GEN_6790; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6792 = 8'h88 == _t_T_50[31:24] ? 8'hc4 : _GEN_6791; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6793 = 8'h89 == _t_T_50[31:24] ? 8'ha7 : _GEN_6792; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6794 = 8'h8a == _t_T_50[31:24] ? 8'h7e : _GEN_6793; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6795 = 8'h8b == _t_T_50[31:24] ? 8'h3d : _GEN_6794; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6796 = 8'h8c == _t_T_50[31:24] ? 8'h64 : _GEN_6795; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6797 = 8'h8d == _t_T_50[31:24] ? 8'h5d : _GEN_6796; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6798 = 8'h8e == _t_T_50[31:24] ? 8'h19 : _GEN_6797; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6799 = 8'h8f == _t_T_50[31:24] ? 8'h73 : _GEN_6798; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6800 = 8'h90 == _t_T_50[31:24] ? 8'h60 : _GEN_6799; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6801 = 8'h91 == _t_T_50[31:24] ? 8'h81 : _GEN_6800; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6802 = 8'h92 == _t_T_50[31:24] ? 8'h4f : _GEN_6801; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6803 = 8'h93 == _t_T_50[31:24] ? 8'hdc : _GEN_6802; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6804 = 8'h94 == _t_T_50[31:24] ? 8'h22 : _GEN_6803; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6805 = 8'h95 == _t_T_50[31:24] ? 8'h2a : _GEN_6804; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6806 = 8'h96 == _t_T_50[31:24] ? 8'h90 : _GEN_6805; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6807 = 8'h97 == _t_T_50[31:24] ? 8'h88 : _GEN_6806; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6808 = 8'h98 == _t_T_50[31:24] ? 8'h46 : _GEN_6807; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6809 = 8'h99 == _t_T_50[31:24] ? 8'hee : _GEN_6808; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6810 = 8'h9a == _t_T_50[31:24] ? 8'hb8 : _GEN_6809; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6811 = 8'h9b == _t_T_50[31:24] ? 8'h14 : _GEN_6810; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6812 = 8'h9c == _t_T_50[31:24] ? 8'hde : _GEN_6811; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6813 = 8'h9d == _t_T_50[31:24] ? 8'h5e : _GEN_6812; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6814 = 8'h9e == _t_T_50[31:24] ? 8'hb : _GEN_6813; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6815 = 8'h9f == _t_T_50[31:24] ? 8'hdb : _GEN_6814; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6816 = 8'ha0 == _t_T_50[31:24] ? 8'he0 : _GEN_6815; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6817 = 8'ha1 == _t_T_50[31:24] ? 8'h32 : _GEN_6816; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6818 = 8'ha2 == _t_T_50[31:24] ? 8'h3a : _GEN_6817; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6819 = 8'ha3 == _t_T_50[31:24] ? 8'ha : _GEN_6818; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6820 = 8'ha4 == _t_T_50[31:24] ? 8'h49 : _GEN_6819; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6821 = 8'ha5 == _t_T_50[31:24] ? 8'h6 : _GEN_6820; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6822 = 8'ha6 == _t_T_50[31:24] ? 8'h24 : _GEN_6821; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6823 = 8'ha7 == _t_T_50[31:24] ? 8'h5c : _GEN_6822; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6824 = 8'ha8 == _t_T_50[31:24] ? 8'hc2 : _GEN_6823; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6825 = 8'ha9 == _t_T_50[31:24] ? 8'hd3 : _GEN_6824; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6826 = 8'haa == _t_T_50[31:24] ? 8'hac : _GEN_6825; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6827 = 8'hab == _t_T_50[31:24] ? 8'h62 : _GEN_6826; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6828 = 8'hac == _t_T_50[31:24] ? 8'h91 : _GEN_6827; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6829 = 8'had == _t_T_50[31:24] ? 8'h95 : _GEN_6828; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6830 = 8'hae == _t_T_50[31:24] ? 8'he4 : _GEN_6829; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6831 = 8'haf == _t_T_50[31:24] ? 8'h79 : _GEN_6830; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6832 = 8'hb0 == _t_T_50[31:24] ? 8'he7 : _GEN_6831; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6833 = 8'hb1 == _t_T_50[31:24] ? 8'hc8 : _GEN_6832; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6834 = 8'hb2 == _t_T_50[31:24] ? 8'h37 : _GEN_6833; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6835 = 8'hb3 == _t_T_50[31:24] ? 8'h6d : _GEN_6834; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6836 = 8'hb4 == _t_T_50[31:24] ? 8'h8d : _GEN_6835; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6837 = 8'hb5 == _t_T_50[31:24] ? 8'hd5 : _GEN_6836; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6838 = 8'hb6 == _t_T_50[31:24] ? 8'h4e : _GEN_6837; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6839 = 8'hb7 == _t_T_50[31:24] ? 8'ha9 : _GEN_6838; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6840 = 8'hb8 == _t_T_50[31:24] ? 8'h6c : _GEN_6839; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6841 = 8'hb9 == _t_T_50[31:24] ? 8'h56 : _GEN_6840; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6842 = 8'hba == _t_T_50[31:24] ? 8'hf4 : _GEN_6841; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6843 = 8'hbb == _t_T_50[31:24] ? 8'hea : _GEN_6842; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6844 = 8'hbc == _t_T_50[31:24] ? 8'h65 : _GEN_6843; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6845 = 8'hbd == _t_T_50[31:24] ? 8'h7a : _GEN_6844; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6846 = 8'hbe == _t_T_50[31:24] ? 8'hae : _GEN_6845; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6847 = 8'hbf == _t_T_50[31:24] ? 8'h8 : _GEN_6846; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6848 = 8'hc0 == _t_T_50[31:24] ? 8'hba : _GEN_6847; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6849 = 8'hc1 == _t_T_50[31:24] ? 8'h78 : _GEN_6848; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6850 = 8'hc2 == _t_T_50[31:24] ? 8'h25 : _GEN_6849; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6851 = 8'hc3 == _t_T_50[31:24] ? 8'h2e : _GEN_6850; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6852 = 8'hc4 == _t_T_50[31:24] ? 8'h1c : _GEN_6851; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6853 = 8'hc5 == _t_T_50[31:24] ? 8'ha6 : _GEN_6852; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6854 = 8'hc6 == _t_T_50[31:24] ? 8'hb4 : _GEN_6853; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6855 = 8'hc7 == _t_T_50[31:24] ? 8'hc6 : _GEN_6854; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6856 = 8'hc8 == _t_T_50[31:24] ? 8'he8 : _GEN_6855; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6857 = 8'hc9 == _t_T_50[31:24] ? 8'hdd : _GEN_6856; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6858 = 8'hca == _t_T_50[31:24] ? 8'h74 : _GEN_6857; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6859 = 8'hcb == _t_T_50[31:24] ? 8'h1f : _GEN_6858; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6860 = 8'hcc == _t_T_50[31:24] ? 8'h4b : _GEN_6859; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6861 = 8'hcd == _t_T_50[31:24] ? 8'hbd : _GEN_6860; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6862 = 8'hce == _t_T_50[31:24] ? 8'h8b : _GEN_6861; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6863 = 8'hcf == _t_T_50[31:24] ? 8'h8a : _GEN_6862; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6864 = 8'hd0 == _t_T_50[31:24] ? 8'h70 : _GEN_6863; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6865 = 8'hd1 == _t_T_50[31:24] ? 8'h3e : _GEN_6864; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6866 = 8'hd2 == _t_T_50[31:24] ? 8'hb5 : _GEN_6865; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6867 = 8'hd3 == _t_T_50[31:24] ? 8'h66 : _GEN_6866; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6868 = 8'hd4 == _t_T_50[31:24] ? 8'h48 : _GEN_6867; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6869 = 8'hd5 == _t_T_50[31:24] ? 8'h3 : _GEN_6868; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6870 = 8'hd6 == _t_T_50[31:24] ? 8'hf6 : _GEN_6869; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6871 = 8'hd7 == _t_T_50[31:24] ? 8'he : _GEN_6870; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6872 = 8'hd8 == _t_T_50[31:24] ? 8'h61 : _GEN_6871; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6873 = 8'hd9 == _t_T_50[31:24] ? 8'h35 : _GEN_6872; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6874 = 8'hda == _t_T_50[31:24] ? 8'h57 : _GEN_6873; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6875 = 8'hdb == _t_T_50[31:24] ? 8'hb9 : _GEN_6874; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6876 = 8'hdc == _t_T_50[31:24] ? 8'h86 : _GEN_6875; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6877 = 8'hdd == _t_T_50[31:24] ? 8'hc1 : _GEN_6876; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6878 = 8'hde == _t_T_50[31:24] ? 8'h1d : _GEN_6877; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6879 = 8'hdf == _t_T_50[31:24] ? 8'h9e : _GEN_6878; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6880 = 8'he0 == _t_T_50[31:24] ? 8'he1 : _GEN_6879; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6881 = 8'he1 == _t_T_50[31:24] ? 8'hf8 : _GEN_6880; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6882 = 8'he2 == _t_T_50[31:24] ? 8'h98 : _GEN_6881; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6883 = 8'he3 == _t_T_50[31:24] ? 8'h11 : _GEN_6882; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6884 = 8'he4 == _t_T_50[31:24] ? 8'h69 : _GEN_6883; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6885 = 8'he5 == _t_T_50[31:24] ? 8'hd9 : _GEN_6884; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6886 = 8'he6 == _t_T_50[31:24] ? 8'h8e : _GEN_6885; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6887 = 8'he7 == _t_T_50[31:24] ? 8'h94 : _GEN_6886; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6888 = 8'he8 == _t_T_50[31:24] ? 8'h9b : _GEN_6887; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6889 = 8'he9 == _t_T_50[31:24] ? 8'h1e : _GEN_6888; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6890 = 8'hea == _t_T_50[31:24] ? 8'h87 : _GEN_6889; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6891 = 8'heb == _t_T_50[31:24] ? 8'he9 : _GEN_6890; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6892 = 8'hec == _t_T_50[31:24] ? 8'hce : _GEN_6891; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6893 = 8'hed == _t_T_50[31:24] ? 8'h55 : _GEN_6892; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6894 = 8'hee == _t_T_50[31:24] ? 8'h28 : _GEN_6893; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6895 = 8'hef == _t_T_50[31:24] ? 8'hdf : _GEN_6894; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6896 = 8'hf0 == _t_T_50[31:24] ? 8'h8c : _GEN_6895; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6897 = 8'hf1 == _t_T_50[31:24] ? 8'ha1 : _GEN_6896; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6898 = 8'hf2 == _t_T_50[31:24] ? 8'h89 : _GEN_6897; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6899 = 8'hf3 == _t_T_50[31:24] ? 8'hd : _GEN_6898; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6900 = 8'hf4 == _t_T_50[31:24] ? 8'hbf : _GEN_6899; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6901 = 8'hf5 == _t_T_50[31:24] ? 8'he6 : _GEN_6900; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6902 = 8'hf6 == _t_T_50[31:24] ? 8'h42 : _GEN_6901; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6903 = 8'hf7 == _t_T_50[31:24] ? 8'h68 : _GEN_6902; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6904 = 8'hf8 == _t_T_50[31:24] ? 8'h41 : _GEN_6903; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6905 = 8'hf9 == _t_T_50[31:24] ? 8'h99 : _GEN_6904; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6906 = 8'hfa == _t_T_50[31:24] ? 8'h2d : _GEN_6905; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6907 = 8'hfb == _t_T_50[31:24] ? 8'hf : _GEN_6906; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6908 = 8'hfc == _t_T_50[31:24] ? 8'hb0 : _GEN_6907; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6909 = 8'hfd == _t_T_50[31:24] ? 8'h54 : _GEN_6908; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6910 = 8'hfe == _t_T_50[31:24] ? 8'hbb : _GEN_6909; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6911 = 8'hff == _t_T_50[31:24] ? 8'h16 : _GEN_6910; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6913 = 8'h1 == _t_T_50[23:16] ? 8'h7c : 8'h63; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6914 = 8'h2 == _t_T_50[23:16] ? 8'h77 : _GEN_6913; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6915 = 8'h3 == _t_T_50[23:16] ? 8'h7b : _GEN_6914; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6916 = 8'h4 == _t_T_50[23:16] ? 8'hf2 : _GEN_6915; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6917 = 8'h5 == _t_T_50[23:16] ? 8'h6b : _GEN_6916; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6918 = 8'h6 == _t_T_50[23:16] ? 8'h6f : _GEN_6917; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6919 = 8'h7 == _t_T_50[23:16] ? 8'hc5 : _GEN_6918; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6920 = 8'h8 == _t_T_50[23:16] ? 8'h30 : _GEN_6919; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6921 = 8'h9 == _t_T_50[23:16] ? 8'h1 : _GEN_6920; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6922 = 8'ha == _t_T_50[23:16] ? 8'h67 : _GEN_6921; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6923 = 8'hb == _t_T_50[23:16] ? 8'h2b : _GEN_6922; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6924 = 8'hc == _t_T_50[23:16] ? 8'hfe : _GEN_6923; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6925 = 8'hd == _t_T_50[23:16] ? 8'hd7 : _GEN_6924; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6926 = 8'he == _t_T_50[23:16] ? 8'hab : _GEN_6925; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6927 = 8'hf == _t_T_50[23:16] ? 8'h76 : _GEN_6926; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6928 = 8'h10 == _t_T_50[23:16] ? 8'hca : _GEN_6927; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6929 = 8'h11 == _t_T_50[23:16] ? 8'h82 : _GEN_6928; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6930 = 8'h12 == _t_T_50[23:16] ? 8'hc9 : _GEN_6929; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6931 = 8'h13 == _t_T_50[23:16] ? 8'h7d : _GEN_6930; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6932 = 8'h14 == _t_T_50[23:16] ? 8'hfa : _GEN_6931; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6933 = 8'h15 == _t_T_50[23:16] ? 8'h59 : _GEN_6932; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6934 = 8'h16 == _t_T_50[23:16] ? 8'h47 : _GEN_6933; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6935 = 8'h17 == _t_T_50[23:16] ? 8'hf0 : _GEN_6934; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6936 = 8'h18 == _t_T_50[23:16] ? 8'had : _GEN_6935; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6937 = 8'h19 == _t_T_50[23:16] ? 8'hd4 : _GEN_6936; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6938 = 8'h1a == _t_T_50[23:16] ? 8'ha2 : _GEN_6937; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6939 = 8'h1b == _t_T_50[23:16] ? 8'haf : _GEN_6938; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6940 = 8'h1c == _t_T_50[23:16] ? 8'h9c : _GEN_6939; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6941 = 8'h1d == _t_T_50[23:16] ? 8'ha4 : _GEN_6940; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6942 = 8'h1e == _t_T_50[23:16] ? 8'h72 : _GEN_6941; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6943 = 8'h1f == _t_T_50[23:16] ? 8'hc0 : _GEN_6942; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6944 = 8'h20 == _t_T_50[23:16] ? 8'hb7 : _GEN_6943; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6945 = 8'h21 == _t_T_50[23:16] ? 8'hfd : _GEN_6944; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6946 = 8'h22 == _t_T_50[23:16] ? 8'h93 : _GEN_6945; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6947 = 8'h23 == _t_T_50[23:16] ? 8'h26 : _GEN_6946; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6948 = 8'h24 == _t_T_50[23:16] ? 8'h36 : _GEN_6947; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6949 = 8'h25 == _t_T_50[23:16] ? 8'h3f : _GEN_6948; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6950 = 8'h26 == _t_T_50[23:16] ? 8'hf7 : _GEN_6949; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6951 = 8'h27 == _t_T_50[23:16] ? 8'hcc : _GEN_6950; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6952 = 8'h28 == _t_T_50[23:16] ? 8'h34 : _GEN_6951; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6953 = 8'h29 == _t_T_50[23:16] ? 8'ha5 : _GEN_6952; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6954 = 8'h2a == _t_T_50[23:16] ? 8'he5 : _GEN_6953; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6955 = 8'h2b == _t_T_50[23:16] ? 8'hf1 : _GEN_6954; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6956 = 8'h2c == _t_T_50[23:16] ? 8'h71 : _GEN_6955; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6957 = 8'h2d == _t_T_50[23:16] ? 8'hd8 : _GEN_6956; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6958 = 8'h2e == _t_T_50[23:16] ? 8'h31 : _GEN_6957; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6959 = 8'h2f == _t_T_50[23:16] ? 8'h15 : _GEN_6958; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6960 = 8'h30 == _t_T_50[23:16] ? 8'h4 : _GEN_6959; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6961 = 8'h31 == _t_T_50[23:16] ? 8'hc7 : _GEN_6960; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6962 = 8'h32 == _t_T_50[23:16] ? 8'h23 : _GEN_6961; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6963 = 8'h33 == _t_T_50[23:16] ? 8'hc3 : _GEN_6962; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6964 = 8'h34 == _t_T_50[23:16] ? 8'h18 : _GEN_6963; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6965 = 8'h35 == _t_T_50[23:16] ? 8'h96 : _GEN_6964; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6966 = 8'h36 == _t_T_50[23:16] ? 8'h5 : _GEN_6965; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6967 = 8'h37 == _t_T_50[23:16] ? 8'h9a : _GEN_6966; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6968 = 8'h38 == _t_T_50[23:16] ? 8'h7 : _GEN_6967; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6969 = 8'h39 == _t_T_50[23:16] ? 8'h12 : _GEN_6968; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6970 = 8'h3a == _t_T_50[23:16] ? 8'h80 : _GEN_6969; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6971 = 8'h3b == _t_T_50[23:16] ? 8'he2 : _GEN_6970; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6972 = 8'h3c == _t_T_50[23:16] ? 8'heb : _GEN_6971; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6973 = 8'h3d == _t_T_50[23:16] ? 8'h27 : _GEN_6972; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6974 = 8'h3e == _t_T_50[23:16] ? 8'hb2 : _GEN_6973; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6975 = 8'h3f == _t_T_50[23:16] ? 8'h75 : _GEN_6974; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6976 = 8'h40 == _t_T_50[23:16] ? 8'h9 : _GEN_6975; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6977 = 8'h41 == _t_T_50[23:16] ? 8'h83 : _GEN_6976; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6978 = 8'h42 == _t_T_50[23:16] ? 8'h2c : _GEN_6977; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6979 = 8'h43 == _t_T_50[23:16] ? 8'h1a : _GEN_6978; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6980 = 8'h44 == _t_T_50[23:16] ? 8'h1b : _GEN_6979; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6981 = 8'h45 == _t_T_50[23:16] ? 8'h6e : _GEN_6980; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6982 = 8'h46 == _t_T_50[23:16] ? 8'h5a : _GEN_6981; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6983 = 8'h47 == _t_T_50[23:16] ? 8'ha0 : _GEN_6982; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6984 = 8'h48 == _t_T_50[23:16] ? 8'h52 : _GEN_6983; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6985 = 8'h49 == _t_T_50[23:16] ? 8'h3b : _GEN_6984; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6986 = 8'h4a == _t_T_50[23:16] ? 8'hd6 : _GEN_6985; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6987 = 8'h4b == _t_T_50[23:16] ? 8'hb3 : _GEN_6986; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6988 = 8'h4c == _t_T_50[23:16] ? 8'h29 : _GEN_6987; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6989 = 8'h4d == _t_T_50[23:16] ? 8'he3 : _GEN_6988; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6990 = 8'h4e == _t_T_50[23:16] ? 8'h2f : _GEN_6989; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6991 = 8'h4f == _t_T_50[23:16] ? 8'h84 : _GEN_6990; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6992 = 8'h50 == _t_T_50[23:16] ? 8'h53 : _GEN_6991; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6993 = 8'h51 == _t_T_50[23:16] ? 8'hd1 : _GEN_6992; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6994 = 8'h52 == _t_T_50[23:16] ? 8'h0 : _GEN_6993; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6995 = 8'h53 == _t_T_50[23:16] ? 8'hed : _GEN_6994; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6996 = 8'h54 == _t_T_50[23:16] ? 8'h20 : _GEN_6995; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6997 = 8'h55 == _t_T_50[23:16] ? 8'hfc : _GEN_6996; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6998 = 8'h56 == _t_T_50[23:16] ? 8'hb1 : _GEN_6997; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_6999 = 8'h57 == _t_T_50[23:16] ? 8'h5b : _GEN_6998; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7000 = 8'h58 == _t_T_50[23:16] ? 8'h6a : _GEN_6999; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7001 = 8'h59 == _t_T_50[23:16] ? 8'hcb : _GEN_7000; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7002 = 8'h5a == _t_T_50[23:16] ? 8'hbe : _GEN_7001; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7003 = 8'h5b == _t_T_50[23:16] ? 8'h39 : _GEN_7002; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7004 = 8'h5c == _t_T_50[23:16] ? 8'h4a : _GEN_7003; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7005 = 8'h5d == _t_T_50[23:16] ? 8'h4c : _GEN_7004; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7006 = 8'h5e == _t_T_50[23:16] ? 8'h58 : _GEN_7005; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7007 = 8'h5f == _t_T_50[23:16] ? 8'hcf : _GEN_7006; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7008 = 8'h60 == _t_T_50[23:16] ? 8'hd0 : _GEN_7007; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7009 = 8'h61 == _t_T_50[23:16] ? 8'hef : _GEN_7008; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7010 = 8'h62 == _t_T_50[23:16] ? 8'haa : _GEN_7009; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7011 = 8'h63 == _t_T_50[23:16] ? 8'hfb : _GEN_7010; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7012 = 8'h64 == _t_T_50[23:16] ? 8'h43 : _GEN_7011; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7013 = 8'h65 == _t_T_50[23:16] ? 8'h4d : _GEN_7012; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7014 = 8'h66 == _t_T_50[23:16] ? 8'h33 : _GEN_7013; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7015 = 8'h67 == _t_T_50[23:16] ? 8'h85 : _GEN_7014; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7016 = 8'h68 == _t_T_50[23:16] ? 8'h45 : _GEN_7015; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7017 = 8'h69 == _t_T_50[23:16] ? 8'hf9 : _GEN_7016; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7018 = 8'h6a == _t_T_50[23:16] ? 8'h2 : _GEN_7017; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7019 = 8'h6b == _t_T_50[23:16] ? 8'h7f : _GEN_7018; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7020 = 8'h6c == _t_T_50[23:16] ? 8'h50 : _GEN_7019; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7021 = 8'h6d == _t_T_50[23:16] ? 8'h3c : _GEN_7020; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7022 = 8'h6e == _t_T_50[23:16] ? 8'h9f : _GEN_7021; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7023 = 8'h6f == _t_T_50[23:16] ? 8'ha8 : _GEN_7022; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7024 = 8'h70 == _t_T_50[23:16] ? 8'h51 : _GEN_7023; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7025 = 8'h71 == _t_T_50[23:16] ? 8'ha3 : _GEN_7024; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7026 = 8'h72 == _t_T_50[23:16] ? 8'h40 : _GEN_7025; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7027 = 8'h73 == _t_T_50[23:16] ? 8'h8f : _GEN_7026; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7028 = 8'h74 == _t_T_50[23:16] ? 8'h92 : _GEN_7027; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7029 = 8'h75 == _t_T_50[23:16] ? 8'h9d : _GEN_7028; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7030 = 8'h76 == _t_T_50[23:16] ? 8'h38 : _GEN_7029; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7031 = 8'h77 == _t_T_50[23:16] ? 8'hf5 : _GEN_7030; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7032 = 8'h78 == _t_T_50[23:16] ? 8'hbc : _GEN_7031; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7033 = 8'h79 == _t_T_50[23:16] ? 8'hb6 : _GEN_7032; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7034 = 8'h7a == _t_T_50[23:16] ? 8'hda : _GEN_7033; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7035 = 8'h7b == _t_T_50[23:16] ? 8'h21 : _GEN_7034; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7036 = 8'h7c == _t_T_50[23:16] ? 8'h10 : _GEN_7035; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7037 = 8'h7d == _t_T_50[23:16] ? 8'hff : _GEN_7036; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7038 = 8'h7e == _t_T_50[23:16] ? 8'hf3 : _GEN_7037; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7039 = 8'h7f == _t_T_50[23:16] ? 8'hd2 : _GEN_7038; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7040 = 8'h80 == _t_T_50[23:16] ? 8'hcd : _GEN_7039; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7041 = 8'h81 == _t_T_50[23:16] ? 8'hc : _GEN_7040; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7042 = 8'h82 == _t_T_50[23:16] ? 8'h13 : _GEN_7041; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7043 = 8'h83 == _t_T_50[23:16] ? 8'hec : _GEN_7042; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7044 = 8'h84 == _t_T_50[23:16] ? 8'h5f : _GEN_7043; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7045 = 8'h85 == _t_T_50[23:16] ? 8'h97 : _GEN_7044; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7046 = 8'h86 == _t_T_50[23:16] ? 8'h44 : _GEN_7045; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7047 = 8'h87 == _t_T_50[23:16] ? 8'h17 : _GEN_7046; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7048 = 8'h88 == _t_T_50[23:16] ? 8'hc4 : _GEN_7047; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7049 = 8'h89 == _t_T_50[23:16] ? 8'ha7 : _GEN_7048; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7050 = 8'h8a == _t_T_50[23:16] ? 8'h7e : _GEN_7049; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7051 = 8'h8b == _t_T_50[23:16] ? 8'h3d : _GEN_7050; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7052 = 8'h8c == _t_T_50[23:16] ? 8'h64 : _GEN_7051; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7053 = 8'h8d == _t_T_50[23:16] ? 8'h5d : _GEN_7052; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7054 = 8'h8e == _t_T_50[23:16] ? 8'h19 : _GEN_7053; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7055 = 8'h8f == _t_T_50[23:16] ? 8'h73 : _GEN_7054; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7056 = 8'h90 == _t_T_50[23:16] ? 8'h60 : _GEN_7055; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7057 = 8'h91 == _t_T_50[23:16] ? 8'h81 : _GEN_7056; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7058 = 8'h92 == _t_T_50[23:16] ? 8'h4f : _GEN_7057; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7059 = 8'h93 == _t_T_50[23:16] ? 8'hdc : _GEN_7058; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7060 = 8'h94 == _t_T_50[23:16] ? 8'h22 : _GEN_7059; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7061 = 8'h95 == _t_T_50[23:16] ? 8'h2a : _GEN_7060; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7062 = 8'h96 == _t_T_50[23:16] ? 8'h90 : _GEN_7061; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7063 = 8'h97 == _t_T_50[23:16] ? 8'h88 : _GEN_7062; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7064 = 8'h98 == _t_T_50[23:16] ? 8'h46 : _GEN_7063; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7065 = 8'h99 == _t_T_50[23:16] ? 8'hee : _GEN_7064; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7066 = 8'h9a == _t_T_50[23:16] ? 8'hb8 : _GEN_7065; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7067 = 8'h9b == _t_T_50[23:16] ? 8'h14 : _GEN_7066; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7068 = 8'h9c == _t_T_50[23:16] ? 8'hde : _GEN_7067; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7069 = 8'h9d == _t_T_50[23:16] ? 8'h5e : _GEN_7068; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7070 = 8'h9e == _t_T_50[23:16] ? 8'hb : _GEN_7069; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7071 = 8'h9f == _t_T_50[23:16] ? 8'hdb : _GEN_7070; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7072 = 8'ha0 == _t_T_50[23:16] ? 8'he0 : _GEN_7071; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7073 = 8'ha1 == _t_T_50[23:16] ? 8'h32 : _GEN_7072; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7074 = 8'ha2 == _t_T_50[23:16] ? 8'h3a : _GEN_7073; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7075 = 8'ha3 == _t_T_50[23:16] ? 8'ha : _GEN_7074; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7076 = 8'ha4 == _t_T_50[23:16] ? 8'h49 : _GEN_7075; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7077 = 8'ha5 == _t_T_50[23:16] ? 8'h6 : _GEN_7076; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7078 = 8'ha6 == _t_T_50[23:16] ? 8'h24 : _GEN_7077; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7079 = 8'ha7 == _t_T_50[23:16] ? 8'h5c : _GEN_7078; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7080 = 8'ha8 == _t_T_50[23:16] ? 8'hc2 : _GEN_7079; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7081 = 8'ha9 == _t_T_50[23:16] ? 8'hd3 : _GEN_7080; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7082 = 8'haa == _t_T_50[23:16] ? 8'hac : _GEN_7081; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7083 = 8'hab == _t_T_50[23:16] ? 8'h62 : _GEN_7082; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7084 = 8'hac == _t_T_50[23:16] ? 8'h91 : _GEN_7083; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7085 = 8'had == _t_T_50[23:16] ? 8'h95 : _GEN_7084; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7086 = 8'hae == _t_T_50[23:16] ? 8'he4 : _GEN_7085; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7087 = 8'haf == _t_T_50[23:16] ? 8'h79 : _GEN_7086; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7088 = 8'hb0 == _t_T_50[23:16] ? 8'he7 : _GEN_7087; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7089 = 8'hb1 == _t_T_50[23:16] ? 8'hc8 : _GEN_7088; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7090 = 8'hb2 == _t_T_50[23:16] ? 8'h37 : _GEN_7089; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7091 = 8'hb3 == _t_T_50[23:16] ? 8'h6d : _GEN_7090; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7092 = 8'hb4 == _t_T_50[23:16] ? 8'h8d : _GEN_7091; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7093 = 8'hb5 == _t_T_50[23:16] ? 8'hd5 : _GEN_7092; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7094 = 8'hb6 == _t_T_50[23:16] ? 8'h4e : _GEN_7093; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7095 = 8'hb7 == _t_T_50[23:16] ? 8'ha9 : _GEN_7094; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7096 = 8'hb8 == _t_T_50[23:16] ? 8'h6c : _GEN_7095; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7097 = 8'hb9 == _t_T_50[23:16] ? 8'h56 : _GEN_7096; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7098 = 8'hba == _t_T_50[23:16] ? 8'hf4 : _GEN_7097; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7099 = 8'hbb == _t_T_50[23:16] ? 8'hea : _GEN_7098; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7100 = 8'hbc == _t_T_50[23:16] ? 8'h65 : _GEN_7099; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7101 = 8'hbd == _t_T_50[23:16] ? 8'h7a : _GEN_7100; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7102 = 8'hbe == _t_T_50[23:16] ? 8'hae : _GEN_7101; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7103 = 8'hbf == _t_T_50[23:16] ? 8'h8 : _GEN_7102; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7104 = 8'hc0 == _t_T_50[23:16] ? 8'hba : _GEN_7103; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7105 = 8'hc1 == _t_T_50[23:16] ? 8'h78 : _GEN_7104; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7106 = 8'hc2 == _t_T_50[23:16] ? 8'h25 : _GEN_7105; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7107 = 8'hc3 == _t_T_50[23:16] ? 8'h2e : _GEN_7106; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7108 = 8'hc4 == _t_T_50[23:16] ? 8'h1c : _GEN_7107; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7109 = 8'hc5 == _t_T_50[23:16] ? 8'ha6 : _GEN_7108; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7110 = 8'hc6 == _t_T_50[23:16] ? 8'hb4 : _GEN_7109; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7111 = 8'hc7 == _t_T_50[23:16] ? 8'hc6 : _GEN_7110; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7112 = 8'hc8 == _t_T_50[23:16] ? 8'he8 : _GEN_7111; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7113 = 8'hc9 == _t_T_50[23:16] ? 8'hdd : _GEN_7112; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7114 = 8'hca == _t_T_50[23:16] ? 8'h74 : _GEN_7113; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7115 = 8'hcb == _t_T_50[23:16] ? 8'h1f : _GEN_7114; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7116 = 8'hcc == _t_T_50[23:16] ? 8'h4b : _GEN_7115; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7117 = 8'hcd == _t_T_50[23:16] ? 8'hbd : _GEN_7116; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7118 = 8'hce == _t_T_50[23:16] ? 8'h8b : _GEN_7117; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7119 = 8'hcf == _t_T_50[23:16] ? 8'h8a : _GEN_7118; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7120 = 8'hd0 == _t_T_50[23:16] ? 8'h70 : _GEN_7119; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7121 = 8'hd1 == _t_T_50[23:16] ? 8'h3e : _GEN_7120; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7122 = 8'hd2 == _t_T_50[23:16] ? 8'hb5 : _GEN_7121; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7123 = 8'hd3 == _t_T_50[23:16] ? 8'h66 : _GEN_7122; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7124 = 8'hd4 == _t_T_50[23:16] ? 8'h48 : _GEN_7123; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7125 = 8'hd5 == _t_T_50[23:16] ? 8'h3 : _GEN_7124; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7126 = 8'hd6 == _t_T_50[23:16] ? 8'hf6 : _GEN_7125; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7127 = 8'hd7 == _t_T_50[23:16] ? 8'he : _GEN_7126; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7128 = 8'hd8 == _t_T_50[23:16] ? 8'h61 : _GEN_7127; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7129 = 8'hd9 == _t_T_50[23:16] ? 8'h35 : _GEN_7128; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7130 = 8'hda == _t_T_50[23:16] ? 8'h57 : _GEN_7129; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7131 = 8'hdb == _t_T_50[23:16] ? 8'hb9 : _GEN_7130; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7132 = 8'hdc == _t_T_50[23:16] ? 8'h86 : _GEN_7131; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7133 = 8'hdd == _t_T_50[23:16] ? 8'hc1 : _GEN_7132; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7134 = 8'hde == _t_T_50[23:16] ? 8'h1d : _GEN_7133; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7135 = 8'hdf == _t_T_50[23:16] ? 8'h9e : _GEN_7134; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7136 = 8'he0 == _t_T_50[23:16] ? 8'he1 : _GEN_7135; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7137 = 8'he1 == _t_T_50[23:16] ? 8'hf8 : _GEN_7136; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7138 = 8'he2 == _t_T_50[23:16] ? 8'h98 : _GEN_7137; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7139 = 8'he3 == _t_T_50[23:16] ? 8'h11 : _GEN_7138; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7140 = 8'he4 == _t_T_50[23:16] ? 8'h69 : _GEN_7139; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7141 = 8'he5 == _t_T_50[23:16] ? 8'hd9 : _GEN_7140; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7142 = 8'he6 == _t_T_50[23:16] ? 8'h8e : _GEN_7141; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7143 = 8'he7 == _t_T_50[23:16] ? 8'h94 : _GEN_7142; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7144 = 8'he8 == _t_T_50[23:16] ? 8'h9b : _GEN_7143; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7145 = 8'he9 == _t_T_50[23:16] ? 8'h1e : _GEN_7144; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7146 = 8'hea == _t_T_50[23:16] ? 8'h87 : _GEN_7145; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7147 = 8'heb == _t_T_50[23:16] ? 8'he9 : _GEN_7146; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7148 = 8'hec == _t_T_50[23:16] ? 8'hce : _GEN_7147; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7149 = 8'hed == _t_T_50[23:16] ? 8'h55 : _GEN_7148; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7150 = 8'hee == _t_T_50[23:16] ? 8'h28 : _GEN_7149; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7151 = 8'hef == _t_T_50[23:16] ? 8'hdf : _GEN_7150; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7152 = 8'hf0 == _t_T_50[23:16] ? 8'h8c : _GEN_7151; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7153 = 8'hf1 == _t_T_50[23:16] ? 8'ha1 : _GEN_7152; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7154 = 8'hf2 == _t_T_50[23:16] ? 8'h89 : _GEN_7153; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7155 = 8'hf3 == _t_T_50[23:16] ? 8'hd : _GEN_7154; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7156 = 8'hf4 == _t_T_50[23:16] ? 8'hbf : _GEN_7155; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7157 = 8'hf5 == _t_T_50[23:16] ? 8'he6 : _GEN_7156; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7158 = 8'hf6 == _t_T_50[23:16] ? 8'h42 : _GEN_7157; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7159 = 8'hf7 == _t_T_50[23:16] ? 8'h68 : _GEN_7158; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7160 = 8'hf8 == _t_T_50[23:16] ? 8'h41 : _GEN_7159; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7161 = 8'hf9 == _t_T_50[23:16] ? 8'h99 : _GEN_7160; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7162 = 8'hfa == _t_T_50[23:16] ? 8'h2d : _GEN_7161; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7163 = 8'hfb == _t_T_50[23:16] ? 8'hf : _GEN_7162; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7164 = 8'hfc == _t_T_50[23:16] ? 8'hb0 : _GEN_7163; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7165 = 8'hfd == _t_T_50[23:16] ? 8'h54 : _GEN_7164; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7166 = 8'hfe == _t_T_50[23:16] ? 8'hbb : _GEN_7165; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7167 = 8'hff == _t_T_50[23:16] ? 8'h16 : _GEN_7166; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [31:0] _t_T_55 = {_GEN_6911,_GEN_7167,_GEN_6399,_GEN_6655}; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:8]
  wire [31:0] t_6 = _t_T_55 ^ 32'h40000000; // @[src/main/scala/crypto/aes/KeySchedule.scala 59:32]
  wire [31:0] w_28 = w_24 ^ t_6; // @[src/main/scala/crypto/aes/KeySchedule.scala 63:21]
  wire [31:0] w_29 = w_25 ^ w_28; // @[src/main/scala/crypto/aes/KeySchedule.scala 63:21]
  wire [31:0] w_30 = w_26 ^ w_29; // @[src/main/scala/crypto/aes/KeySchedule.scala 63:21]
  wire [31:0] w_31 = w_27 ^ w_30; // @[src/main/scala/crypto/aes/KeySchedule.scala 63:21]
  wire [31:0] _t_T_58 = {w_31[23:0],w_31[31:24]}; // @[src/main/scala/crypto/aes/KeySchedule.scala 23:43]
  wire [7:0] _GEN_7169 = 8'h1 == _t_T_58[15:8] ? 8'h7c : 8'h63; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7170 = 8'h2 == _t_T_58[15:8] ? 8'h77 : _GEN_7169; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7171 = 8'h3 == _t_T_58[15:8] ? 8'h7b : _GEN_7170; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7172 = 8'h4 == _t_T_58[15:8] ? 8'hf2 : _GEN_7171; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7173 = 8'h5 == _t_T_58[15:8] ? 8'h6b : _GEN_7172; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7174 = 8'h6 == _t_T_58[15:8] ? 8'h6f : _GEN_7173; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7175 = 8'h7 == _t_T_58[15:8] ? 8'hc5 : _GEN_7174; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7176 = 8'h8 == _t_T_58[15:8] ? 8'h30 : _GEN_7175; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7177 = 8'h9 == _t_T_58[15:8] ? 8'h1 : _GEN_7176; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7178 = 8'ha == _t_T_58[15:8] ? 8'h67 : _GEN_7177; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7179 = 8'hb == _t_T_58[15:8] ? 8'h2b : _GEN_7178; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7180 = 8'hc == _t_T_58[15:8] ? 8'hfe : _GEN_7179; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7181 = 8'hd == _t_T_58[15:8] ? 8'hd7 : _GEN_7180; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7182 = 8'he == _t_T_58[15:8] ? 8'hab : _GEN_7181; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7183 = 8'hf == _t_T_58[15:8] ? 8'h76 : _GEN_7182; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7184 = 8'h10 == _t_T_58[15:8] ? 8'hca : _GEN_7183; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7185 = 8'h11 == _t_T_58[15:8] ? 8'h82 : _GEN_7184; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7186 = 8'h12 == _t_T_58[15:8] ? 8'hc9 : _GEN_7185; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7187 = 8'h13 == _t_T_58[15:8] ? 8'h7d : _GEN_7186; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7188 = 8'h14 == _t_T_58[15:8] ? 8'hfa : _GEN_7187; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7189 = 8'h15 == _t_T_58[15:8] ? 8'h59 : _GEN_7188; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7190 = 8'h16 == _t_T_58[15:8] ? 8'h47 : _GEN_7189; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7191 = 8'h17 == _t_T_58[15:8] ? 8'hf0 : _GEN_7190; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7192 = 8'h18 == _t_T_58[15:8] ? 8'had : _GEN_7191; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7193 = 8'h19 == _t_T_58[15:8] ? 8'hd4 : _GEN_7192; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7194 = 8'h1a == _t_T_58[15:8] ? 8'ha2 : _GEN_7193; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7195 = 8'h1b == _t_T_58[15:8] ? 8'haf : _GEN_7194; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7196 = 8'h1c == _t_T_58[15:8] ? 8'h9c : _GEN_7195; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7197 = 8'h1d == _t_T_58[15:8] ? 8'ha4 : _GEN_7196; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7198 = 8'h1e == _t_T_58[15:8] ? 8'h72 : _GEN_7197; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7199 = 8'h1f == _t_T_58[15:8] ? 8'hc0 : _GEN_7198; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7200 = 8'h20 == _t_T_58[15:8] ? 8'hb7 : _GEN_7199; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7201 = 8'h21 == _t_T_58[15:8] ? 8'hfd : _GEN_7200; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7202 = 8'h22 == _t_T_58[15:8] ? 8'h93 : _GEN_7201; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7203 = 8'h23 == _t_T_58[15:8] ? 8'h26 : _GEN_7202; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7204 = 8'h24 == _t_T_58[15:8] ? 8'h36 : _GEN_7203; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7205 = 8'h25 == _t_T_58[15:8] ? 8'h3f : _GEN_7204; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7206 = 8'h26 == _t_T_58[15:8] ? 8'hf7 : _GEN_7205; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7207 = 8'h27 == _t_T_58[15:8] ? 8'hcc : _GEN_7206; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7208 = 8'h28 == _t_T_58[15:8] ? 8'h34 : _GEN_7207; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7209 = 8'h29 == _t_T_58[15:8] ? 8'ha5 : _GEN_7208; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7210 = 8'h2a == _t_T_58[15:8] ? 8'he5 : _GEN_7209; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7211 = 8'h2b == _t_T_58[15:8] ? 8'hf1 : _GEN_7210; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7212 = 8'h2c == _t_T_58[15:8] ? 8'h71 : _GEN_7211; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7213 = 8'h2d == _t_T_58[15:8] ? 8'hd8 : _GEN_7212; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7214 = 8'h2e == _t_T_58[15:8] ? 8'h31 : _GEN_7213; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7215 = 8'h2f == _t_T_58[15:8] ? 8'h15 : _GEN_7214; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7216 = 8'h30 == _t_T_58[15:8] ? 8'h4 : _GEN_7215; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7217 = 8'h31 == _t_T_58[15:8] ? 8'hc7 : _GEN_7216; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7218 = 8'h32 == _t_T_58[15:8] ? 8'h23 : _GEN_7217; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7219 = 8'h33 == _t_T_58[15:8] ? 8'hc3 : _GEN_7218; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7220 = 8'h34 == _t_T_58[15:8] ? 8'h18 : _GEN_7219; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7221 = 8'h35 == _t_T_58[15:8] ? 8'h96 : _GEN_7220; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7222 = 8'h36 == _t_T_58[15:8] ? 8'h5 : _GEN_7221; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7223 = 8'h37 == _t_T_58[15:8] ? 8'h9a : _GEN_7222; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7224 = 8'h38 == _t_T_58[15:8] ? 8'h7 : _GEN_7223; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7225 = 8'h39 == _t_T_58[15:8] ? 8'h12 : _GEN_7224; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7226 = 8'h3a == _t_T_58[15:8] ? 8'h80 : _GEN_7225; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7227 = 8'h3b == _t_T_58[15:8] ? 8'he2 : _GEN_7226; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7228 = 8'h3c == _t_T_58[15:8] ? 8'heb : _GEN_7227; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7229 = 8'h3d == _t_T_58[15:8] ? 8'h27 : _GEN_7228; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7230 = 8'h3e == _t_T_58[15:8] ? 8'hb2 : _GEN_7229; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7231 = 8'h3f == _t_T_58[15:8] ? 8'h75 : _GEN_7230; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7232 = 8'h40 == _t_T_58[15:8] ? 8'h9 : _GEN_7231; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7233 = 8'h41 == _t_T_58[15:8] ? 8'h83 : _GEN_7232; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7234 = 8'h42 == _t_T_58[15:8] ? 8'h2c : _GEN_7233; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7235 = 8'h43 == _t_T_58[15:8] ? 8'h1a : _GEN_7234; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7236 = 8'h44 == _t_T_58[15:8] ? 8'h1b : _GEN_7235; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7237 = 8'h45 == _t_T_58[15:8] ? 8'h6e : _GEN_7236; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7238 = 8'h46 == _t_T_58[15:8] ? 8'h5a : _GEN_7237; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7239 = 8'h47 == _t_T_58[15:8] ? 8'ha0 : _GEN_7238; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7240 = 8'h48 == _t_T_58[15:8] ? 8'h52 : _GEN_7239; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7241 = 8'h49 == _t_T_58[15:8] ? 8'h3b : _GEN_7240; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7242 = 8'h4a == _t_T_58[15:8] ? 8'hd6 : _GEN_7241; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7243 = 8'h4b == _t_T_58[15:8] ? 8'hb3 : _GEN_7242; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7244 = 8'h4c == _t_T_58[15:8] ? 8'h29 : _GEN_7243; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7245 = 8'h4d == _t_T_58[15:8] ? 8'he3 : _GEN_7244; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7246 = 8'h4e == _t_T_58[15:8] ? 8'h2f : _GEN_7245; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7247 = 8'h4f == _t_T_58[15:8] ? 8'h84 : _GEN_7246; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7248 = 8'h50 == _t_T_58[15:8] ? 8'h53 : _GEN_7247; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7249 = 8'h51 == _t_T_58[15:8] ? 8'hd1 : _GEN_7248; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7250 = 8'h52 == _t_T_58[15:8] ? 8'h0 : _GEN_7249; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7251 = 8'h53 == _t_T_58[15:8] ? 8'hed : _GEN_7250; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7252 = 8'h54 == _t_T_58[15:8] ? 8'h20 : _GEN_7251; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7253 = 8'h55 == _t_T_58[15:8] ? 8'hfc : _GEN_7252; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7254 = 8'h56 == _t_T_58[15:8] ? 8'hb1 : _GEN_7253; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7255 = 8'h57 == _t_T_58[15:8] ? 8'h5b : _GEN_7254; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7256 = 8'h58 == _t_T_58[15:8] ? 8'h6a : _GEN_7255; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7257 = 8'h59 == _t_T_58[15:8] ? 8'hcb : _GEN_7256; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7258 = 8'h5a == _t_T_58[15:8] ? 8'hbe : _GEN_7257; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7259 = 8'h5b == _t_T_58[15:8] ? 8'h39 : _GEN_7258; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7260 = 8'h5c == _t_T_58[15:8] ? 8'h4a : _GEN_7259; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7261 = 8'h5d == _t_T_58[15:8] ? 8'h4c : _GEN_7260; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7262 = 8'h5e == _t_T_58[15:8] ? 8'h58 : _GEN_7261; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7263 = 8'h5f == _t_T_58[15:8] ? 8'hcf : _GEN_7262; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7264 = 8'h60 == _t_T_58[15:8] ? 8'hd0 : _GEN_7263; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7265 = 8'h61 == _t_T_58[15:8] ? 8'hef : _GEN_7264; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7266 = 8'h62 == _t_T_58[15:8] ? 8'haa : _GEN_7265; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7267 = 8'h63 == _t_T_58[15:8] ? 8'hfb : _GEN_7266; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7268 = 8'h64 == _t_T_58[15:8] ? 8'h43 : _GEN_7267; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7269 = 8'h65 == _t_T_58[15:8] ? 8'h4d : _GEN_7268; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7270 = 8'h66 == _t_T_58[15:8] ? 8'h33 : _GEN_7269; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7271 = 8'h67 == _t_T_58[15:8] ? 8'h85 : _GEN_7270; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7272 = 8'h68 == _t_T_58[15:8] ? 8'h45 : _GEN_7271; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7273 = 8'h69 == _t_T_58[15:8] ? 8'hf9 : _GEN_7272; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7274 = 8'h6a == _t_T_58[15:8] ? 8'h2 : _GEN_7273; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7275 = 8'h6b == _t_T_58[15:8] ? 8'h7f : _GEN_7274; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7276 = 8'h6c == _t_T_58[15:8] ? 8'h50 : _GEN_7275; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7277 = 8'h6d == _t_T_58[15:8] ? 8'h3c : _GEN_7276; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7278 = 8'h6e == _t_T_58[15:8] ? 8'h9f : _GEN_7277; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7279 = 8'h6f == _t_T_58[15:8] ? 8'ha8 : _GEN_7278; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7280 = 8'h70 == _t_T_58[15:8] ? 8'h51 : _GEN_7279; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7281 = 8'h71 == _t_T_58[15:8] ? 8'ha3 : _GEN_7280; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7282 = 8'h72 == _t_T_58[15:8] ? 8'h40 : _GEN_7281; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7283 = 8'h73 == _t_T_58[15:8] ? 8'h8f : _GEN_7282; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7284 = 8'h74 == _t_T_58[15:8] ? 8'h92 : _GEN_7283; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7285 = 8'h75 == _t_T_58[15:8] ? 8'h9d : _GEN_7284; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7286 = 8'h76 == _t_T_58[15:8] ? 8'h38 : _GEN_7285; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7287 = 8'h77 == _t_T_58[15:8] ? 8'hf5 : _GEN_7286; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7288 = 8'h78 == _t_T_58[15:8] ? 8'hbc : _GEN_7287; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7289 = 8'h79 == _t_T_58[15:8] ? 8'hb6 : _GEN_7288; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7290 = 8'h7a == _t_T_58[15:8] ? 8'hda : _GEN_7289; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7291 = 8'h7b == _t_T_58[15:8] ? 8'h21 : _GEN_7290; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7292 = 8'h7c == _t_T_58[15:8] ? 8'h10 : _GEN_7291; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7293 = 8'h7d == _t_T_58[15:8] ? 8'hff : _GEN_7292; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7294 = 8'h7e == _t_T_58[15:8] ? 8'hf3 : _GEN_7293; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7295 = 8'h7f == _t_T_58[15:8] ? 8'hd2 : _GEN_7294; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7296 = 8'h80 == _t_T_58[15:8] ? 8'hcd : _GEN_7295; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7297 = 8'h81 == _t_T_58[15:8] ? 8'hc : _GEN_7296; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7298 = 8'h82 == _t_T_58[15:8] ? 8'h13 : _GEN_7297; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7299 = 8'h83 == _t_T_58[15:8] ? 8'hec : _GEN_7298; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7300 = 8'h84 == _t_T_58[15:8] ? 8'h5f : _GEN_7299; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7301 = 8'h85 == _t_T_58[15:8] ? 8'h97 : _GEN_7300; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7302 = 8'h86 == _t_T_58[15:8] ? 8'h44 : _GEN_7301; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7303 = 8'h87 == _t_T_58[15:8] ? 8'h17 : _GEN_7302; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7304 = 8'h88 == _t_T_58[15:8] ? 8'hc4 : _GEN_7303; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7305 = 8'h89 == _t_T_58[15:8] ? 8'ha7 : _GEN_7304; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7306 = 8'h8a == _t_T_58[15:8] ? 8'h7e : _GEN_7305; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7307 = 8'h8b == _t_T_58[15:8] ? 8'h3d : _GEN_7306; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7308 = 8'h8c == _t_T_58[15:8] ? 8'h64 : _GEN_7307; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7309 = 8'h8d == _t_T_58[15:8] ? 8'h5d : _GEN_7308; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7310 = 8'h8e == _t_T_58[15:8] ? 8'h19 : _GEN_7309; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7311 = 8'h8f == _t_T_58[15:8] ? 8'h73 : _GEN_7310; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7312 = 8'h90 == _t_T_58[15:8] ? 8'h60 : _GEN_7311; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7313 = 8'h91 == _t_T_58[15:8] ? 8'h81 : _GEN_7312; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7314 = 8'h92 == _t_T_58[15:8] ? 8'h4f : _GEN_7313; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7315 = 8'h93 == _t_T_58[15:8] ? 8'hdc : _GEN_7314; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7316 = 8'h94 == _t_T_58[15:8] ? 8'h22 : _GEN_7315; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7317 = 8'h95 == _t_T_58[15:8] ? 8'h2a : _GEN_7316; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7318 = 8'h96 == _t_T_58[15:8] ? 8'h90 : _GEN_7317; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7319 = 8'h97 == _t_T_58[15:8] ? 8'h88 : _GEN_7318; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7320 = 8'h98 == _t_T_58[15:8] ? 8'h46 : _GEN_7319; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7321 = 8'h99 == _t_T_58[15:8] ? 8'hee : _GEN_7320; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7322 = 8'h9a == _t_T_58[15:8] ? 8'hb8 : _GEN_7321; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7323 = 8'h9b == _t_T_58[15:8] ? 8'h14 : _GEN_7322; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7324 = 8'h9c == _t_T_58[15:8] ? 8'hde : _GEN_7323; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7325 = 8'h9d == _t_T_58[15:8] ? 8'h5e : _GEN_7324; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7326 = 8'h9e == _t_T_58[15:8] ? 8'hb : _GEN_7325; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7327 = 8'h9f == _t_T_58[15:8] ? 8'hdb : _GEN_7326; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7328 = 8'ha0 == _t_T_58[15:8] ? 8'he0 : _GEN_7327; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7329 = 8'ha1 == _t_T_58[15:8] ? 8'h32 : _GEN_7328; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7330 = 8'ha2 == _t_T_58[15:8] ? 8'h3a : _GEN_7329; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7331 = 8'ha3 == _t_T_58[15:8] ? 8'ha : _GEN_7330; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7332 = 8'ha4 == _t_T_58[15:8] ? 8'h49 : _GEN_7331; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7333 = 8'ha5 == _t_T_58[15:8] ? 8'h6 : _GEN_7332; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7334 = 8'ha6 == _t_T_58[15:8] ? 8'h24 : _GEN_7333; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7335 = 8'ha7 == _t_T_58[15:8] ? 8'h5c : _GEN_7334; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7336 = 8'ha8 == _t_T_58[15:8] ? 8'hc2 : _GEN_7335; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7337 = 8'ha9 == _t_T_58[15:8] ? 8'hd3 : _GEN_7336; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7338 = 8'haa == _t_T_58[15:8] ? 8'hac : _GEN_7337; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7339 = 8'hab == _t_T_58[15:8] ? 8'h62 : _GEN_7338; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7340 = 8'hac == _t_T_58[15:8] ? 8'h91 : _GEN_7339; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7341 = 8'had == _t_T_58[15:8] ? 8'h95 : _GEN_7340; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7342 = 8'hae == _t_T_58[15:8] ? 8'he4 : _GEN_7341; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7343 = 8'haf == _t_T_58[15:8] ? 8'h79 : _GEN_7342; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7344 = 8'hb0 == _t_T_58[15:8] ? 8'he7 : _GEN_7343; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7345 = 8'hb1 == _t_T_58[15:8] ? 8'hc8 : _GEN_7344; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7346 = 8'hb2 == _t_T_58[15:8] ? 8'h37 : _GEN_7345; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7347 = 8'hb3 == _t_T_58[15:8] ? 8'h6d : _GEN_7346; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7348 = 8'hb4 == _t_T_58[15:8] ? 8'h8d : _GEN_7347; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7349 = 8'hb5 == _t_T_58[15:8] ? 8'hd5 : _GEN_7348; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7350 = 8'hb6 == _t_T_58[15:8] ? 8'h4e : _GEN_7349; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7351 = 8'hb7 == _t_T_58[15:8] ? 8'ha9 : _GEN_7350; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7352 = 8'hb8 == _t_T_58[15:8] ? 8'h6c : _GEN_7351; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7353 = 8'hb9 == _t_T_58[15:8] ? 8'h56 : _GEN_7352; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7354 = 8'hba == _t_T_58[15:8] ? 8'hf4 : _GEN_7353; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7355 = 8'hbb == _t_T_58[15:8] ? 8'hea : _GEN_7354; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7356 = 8'hbc == _t_T_58[15:8] ? 8'h65 : _GEN_7355; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7357 = 8'hbd == _t_T_58[15:8] ? 8'h7a : _GEN_7356; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7358 = 8'hbe == _t_T_58[15:8] ? 8'hae : _GEN_7357; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7359 = 8'hbf == _t_T_58[15:8] ? 8'h8 : _GEN_7358; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7360 = 8'hc0 == _t_T_58[15:8] ? 8'hba : _GEN_7359; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7361 = 8'hc1 == _t_T_58[15:8] ? 8'h78 : _GEN_7360; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7362 = 8'hc2 == _t_T_58[15:8] ? 8'h25 : _GEN_7361; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7363 = 8'hc3 == _t_T_58[15:8] ? 8'h2e : _GEN_7362; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7364 = 8'hc4 == _t_T_58[15:8] ? 8'h1c : _GEN_7363; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7365 = 8'hc5 == _t_T_58[15:8] ? 8'ha6 : _GEN_7364; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7366 = 8'hc6 == _t_T_58[15:8] ? 8'hb4 : _GEN_7365; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7367 = 8'hc7 == _t_T_58[15:8] ? 8'hc6 : _GEN_7366; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7368 = 8'hc8 == _t_T_58[15:8] ? 8'he8 : _GEN_7367; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7369 = 8'hc9 == _t_T_58[15:8] ? 8'hdd : _GEN_7368; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7370 = 8'hca == _t_T_58[15:8] ? 8'h74 : _GEN_7369; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7371 = 8'hcb == _t_T_58[15:8] ? 8'h1f : _GEN_7370; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7372 = 8'hcc == _t_T_58[15:8] ? 8'h4b : _GEN_7371; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7373 = 8'hcd == _t_T_58[15:8] ? 8'hbd : _GEN_7372; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7374 = 8'hce == _t_T_58[15:8] ? 8'h8b : _GEN_7373; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7375 = 8'hcf == _t_T_58[15:8] ? 8'h8a : _GEN_7374; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7376 = 8'hd0 == _t_T_58[15:8] ? 8'h70 : _GEN_7375; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7377 = 8'hd1 == _t_T_58[15:8] ? 8'h3e : _GEN_7376; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7378 = 8'hd2 == _t_T_58[15:8] ? 8'hb5 : _GEN_7377; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7379 = 8'hd3 == _t_T_58[15:8] ? 8'h66 : _GEN_7378; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7380 = 8'hd4 == _t_T_58[15:8] ? 8'h48 : _GEN_7379; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7381 = 8'hd5 == _t_T_58[15:8] ? 8'h3 : _GEN_7380; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7382 = 8'hd6 == _t_T_58[15:8] ? 8'hf6 : _GEN_7381; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7383 = 8'hd7 == _t_T_58[15:8] ? 8'he : _GEN_7382; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7384 = 8'hd8 == _t_T_58[15:8] ? 8'h61 : _GEN_7383; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7385 = 8'hd9 == _t_T_58[15:8] ? 8'h35 : _GEN_7384; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7386 = 8'hda == _t_T_58[15:8] ? 8'h57 : _GEN_7385; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7387 = 8'hdb == _t_T_58[15:8] ? 8'hb9 : _GEN_7386; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7388 = 8'hdc == _t_T_58[15:8] ? 8'h86 : _GEN_7387; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7389 = 8'hdd == _t_T_58[15:8] ? 8'hc1 : _GEN_7388; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7390 = 8'hde == _t_T_58[15:8] ? 8'h1d : _GEN_7389; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7391 = 8'hdf == _t_T_58[15:8] ? 8'h9e : _GEN_7390; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7392 = 8'he0 == _t_T_58[15:8] ? 8'he1 : _GEN_7391; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7393 = 8'he1 == _t_T_58[15:8] ? 8'hf8 : _GEN_7392; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7394 = 8'he2 == _t_T_58[15:8] ? 8'h98 : _GEN_7393; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7395 = 8'he3 == _t_T_58[15:8] ? 8'h11 : _GEN_7394; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7396 = 8'he4 == _t_T_58[15:8] ? 8'h69 : _GEN_7395; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7397 = 8'he5 == _t_T_58[15:8] ? 8'hd9 : _GEN_7396; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7398 = 8'he6 == _t_T_58[15:8] ? 8'h8e : _GEN_7397; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7399 = 8'he7 == _t_T_58[15:8] ? 8'h94 : _GEN_7398; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7400 = 8'he8 == _t_T_58[15:8] ? 8'h9b : _GEN_7399; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7401 = 8'he9 == _t_T_58[15:8] ? 8'h1e : _GEN_7400; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7402 = 8'hea == _t_T_58[15:8] ? 8'h87 : _GEN_7401; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7403 = 8'heb == _t_T_58[15:8] ? 8'he9 : _GEN_7402; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7404 = 8'hec == _t_T_58[15:8] ? 8'hce : _GEN_7403; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7405 = 8'hed == _t_T_58[15:8] ? 8'h55 : _GEN_7404; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7406 = 8'hee == _t_T_58[15:8] ? 8'h28 : _GEN_7405; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7407 = 8'hef == _t_T_58[15:8] ? 8'hdf : _GEN_7406; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7408 = 8'hf0 == _t_T_58[15:8] ? 8'h8c : _GEN_7407; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7409 = 8'hf1 == _t_T_58[15:8] ? 8'ha1 : _GEN_7408; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7410 = 8'hf2 == _t_T_58[15:8] ? 8'h89 : _GEN_7409; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7411 = 8'hf3 == _t_T_58[15:8] ? 8'hd : _GEN_7410; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7412 = 8'hf4 == _t_T_58[15:8] ? 8'hbf : _GEN_7411; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7413 = 8'hf5 == _t_T_58[15:8] ? 8'he6 : _GEN_7412; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7414 = 8'hf6 == _t_T_58[15:8] ? 8'h42 : _GEN_7413; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7415 = 8'hf7 == _t_T_58[15:8] ? 8'h68 : _GEN_7414; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7416 = 8'hf8 == _t_T_58[15:8] ? 8'h41 : _GEN_7415; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7417 = 8'hf9 == _t_T_58[15:8] ? 8'h99 : _GEN_7416; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7418 = 8'hfa == _t_T_58[15:8] ? 8'h2d : _GEN_7417; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7419 = 8'hfb == _t_T_58[15:8] ? 8'hf : _GEN_7418; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7420 = 8'hfc == _t_T_58[15:8] ? 8'hb0 : _GEN_7419; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7421 = 8'hfd == _t_T_58[15:8] ? 8'h54 : _GEN_7420; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7422 = 8'hfe == _t_T_58[15:8] ? 8'hbb : _GEN_7421; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7423 = 8'hff == _t_T_58[15:8] ? 8'h16 : _GEN_7422; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7425 = 8'h1 == _t_T_58[7:0] ? 8'h7c : 8'h63; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7426 = 8'h2 == _t_T_58[7:0] ? 8'h77 : _GEN_7425; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7427 = 8'h3 == _t_T_58[7:0] ? 8'h7b : _GEN_7426; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7428 = 8'h4 == _t_T_58[7:0] ? 8'hf2 : _GEN_7427; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7429 = 8'h5 == _t_T_58[7:0] ? 8'h6b : _GEN_7428; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7430 = 8'h6 == _t_T_58[7:0] ? 8'h6f : _GEN_7429; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7431 = 8'h7 == _t_T_58[7:0] ? 8'hc5 : _GEN_7430; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7432 = 8'h8 == _t_T_58[7:0] ? 8'h30 : _GEN_7431; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7433 = 8'h9 == _t_T_58[7:0] ? 8'h1 : _GEN_7432; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7434 = 8'ha == _t_T_58[7:0] ? 8'h67 : _GEN_7433; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7435 = 8'hb == _t_T_58[7:0] ? 8'h2b : _GEN_7434; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7436 = 8'hc == _t_T_58[7:0] ? 8'hfe : _GEN_7435; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7437 = 8'hd == _t_T_58[7:0] ? 8'hd7 : _GEN_7436; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7438 = 8'he == _t_T_58[7:0] ? 8'hab : _GEN_7437; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7439 = 8'hf == _t_T_58[7:0] ? 8'h76 : _GEN_7438; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7440 = 8'h10 == _t_T_58[7:0] ? 8'hca : _GEN_7439; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7441 = 8'h11 == _t_T_58[7:0] ? 8'h82 : _GEN_7440; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7442 = 8'h12 == _t_T_58[7:0] ? 8'hc9 : _GEN_7441; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7443 = 8'h13 == _t_T_58[7:0] ? 8'h7d : _GEN_7442; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7444 = 8'h14 == _t_T_58[7:0] ? 8'hfa : _GEN_7443; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7445 = 8'h15 == _t_T_58[7:0] ? 8'h59 : _GEN_7444; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7446 = 8'h16 == _t_T_58[7:0] ? 8'h47 : _GEN_7445; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7447 = 8'h17 == _t_T_58[7:0] ? 8'hf0 : _GEN_7446; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7448 = 8'h18 == _t_T_58[7:0] ? 8'had : _GEN_7447; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7449 = 8'h19 == _t_T_58[7:0] ? 8'hd4 : _GEN_7448; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7450 = 8'h1a == _t_T_58[7:0] ? 8'ha2 : _GEN_7449; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7451 = 8'h1b == _t_T_58[7:0] ? 8'haf : _GEN_7450; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7452 = 8'h1c == _t_T_58[7:0] ? 8'h9c : _GEN_7451; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7453 = 8'h1d == _t_T_58[7:0] ? 8'ha4 : _GEN_7452; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7454 = 8'h1e == _t_T_58[7:0] ? 8'h72 : _GEN_7453; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7455 = 8'h1f == _t_T_58[7:0] ? 8'hc0 : _GEN_7454; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7456 = 8'h20 == _t_T_58[7:0] ? 8'hb7 : _GEN_7455; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7457 = 8'h21 == _t_T_58[7:0] ? 8'hfd : _GEN_7456; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7458 = 8'h22 == _t_T_58[7:0] ? 8'h93 : _GEN_7457; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7459 = 8'h23 == _t_T_58[7:0] ? 8'h26 : _GEN_7458; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7460 = 8'h24 == _t_T_58[7:0] ? 8'h36 : _GEN_7459; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7461 = 8'h25 == _t_T_58[7:0] ? 8'h3f : _GEN_7460; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7462 = 8'h26 == _t_T_58[7:0] ? 8'hf7 : _GEN_7461; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7463 = 8'h27 == _t_T_58[7:0] ? 8'hcc : _GEN_7462; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7464 = 8'h28 == _t_T_58[7:0] ? 8'h34 : _GEN_7463; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7465 = 8'h29 == _t_T_58[7:0] ? 8'ha5 : _GEN_7464; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7466 = 8'h2a == _t_T_58[7:0] ? 8'he5 : _GEN_7465; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7467 = 8'h2b == _t_T_58[7:0] ? 8'hf1 : _GEN_7466; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7468 = 8'h2c == _t_T_58[7:0] ? 8'h71 : _GEN_7467; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7469 = 8'h2d == _t_T_58[7:0] ? 8'hd8 : _GEN_7468; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7470 = 8'h2e == _t_T_58[7:0] ? 8'h31 : _GEN_7469; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7471 = 8'h2f == _t_T_58[7:0] ? 8'h15 : _GEN_7470; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7472 = 8'h30 == _t_T_58[7:0] ? 8'h4 : _GEN_7471; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7473 = 8'h31 == _t_T_58[7:0] ? 8'hc7 : _GEN_7472; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7474 = 8'h32 == _t_T_58[7:0] ? 8'h23 : _GEN_7473; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7475 = 8'h33 == _t_T_58[7:0] ? 8'hc3 : _GEN_7474; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7476 = 8'h34 == _t_T_58[7:0] ? 8'h18 : _GEN_7475; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7477 = 8'h35 == _t_T_58[7:0] ? 8'h96 : _GEN_7476; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7478 = 8'h36 == _t_T_58[7:0] ? 8'h5 : _GEN_7477; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7479 = 8'h37 == _t_T_58[7:0] ? 8'h9a : _GEN_7478; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7480 = 8'h38 == _t_T_58[7:0] ? 8'h7 : _GEN_7479; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7481 = 8'h39 == _t_T_58[7:0] ? 8'h12 : _GEN_7480; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7482 = 8'h3a == _t_T_58[7:0] ? 8'h80 : _GEN_7481; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7483 = 8'h3b == _t_T_58[7:0] ? 8'he2 : _GEN_7482; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7484 = 8'h3c == _t_T_58[7:0] ? 8'heb : _GEN_7483; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7485 = 8'h3d == _t_T_58[7:0] ? 8'h27 : _GEN_7484; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7486 = 8'h3e == _t_T_58[7:0] ? 8'hb2 : _GEN_7485; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7487 = 8'h3f == _t_T_58[7:0] ? 8'h75 : _GEN_7486; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7488 = 8'h40 == _t_T_58[7:0] ? 8'h9 : _GEN_7487; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7489 = 8'h41 == _t_T_58[7:0] ? 8'h83 : _GEN_7488; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7490 = 8'h42 == _t_T_58[7:0] ? 8'h2c : _GEN_7489; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7491 = 8'h43 == _t_T_58[7:0] ? 8'h1a : _GEN_7490; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7492 = 8'h44 == _t_T_58[7:0] ? 8'h1b : _GEN_7491; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7493 = 8'h45 == _t_T_58[7:0] ? 8'h6e : _GEN_7492; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7494 = 8'h46 == _t_T_58[7:0] ? 8'h5a : _GEN_7493; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7495 = 8'h47 == _t_T_58[7:0] ? 8'ha0 : _GEN_7494; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7496 = 8'h48 == _t_T_58[7:0] ? 8'h52 : _GEN_7495; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7497 = 8'h49 == _t_T_58[7:0] ? 8'h3b : _GEN_7496; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7498 = 8'h4a == _t_T_58[7:0] ? 8'hd6 : _GEN_7497; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7499 = 8'h4b == _t_T_58[7:0] ? 8'hb3 : _GEN_7498; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7500 = 8'h4c == _t_T_58[7:0] ? 8'h29 : _GEN_7499; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7501 = 8'h4d == _t_T_58[7:0] ? 8'he3 : _GEN_7500; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7502 = 8'h4e == _t_T_58[7:0] ? 8'h2f : _GEN_7501; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7503 = 8'h4f == _t_T_58[7:0] ? 8'h84 : _GEN_7502; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7504 = 8'h50 == _t_T_58[7:0] ? 8'h53 : _GEN_7503; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7505 = 8'h51 == _t_T_58[7:0] ? 8'hd1 : _GEN_7504; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7506 = 8'h52 == _t_T_58[7:0] ? 8'h0 : _GEN_7505; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7507 = 8'h53 == _t_T_58[7:0] ? 8'hed : _GEN_7506; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7508 = 8'h54 == _t_T_58[7:0] ? 8'h20 : _GEN_7507; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7509 = 8'h55 == _t_T_58[7:0] ? 8'hfc : _GEN_7508; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7510 = 8'h56 == _t_T_58[7:0] ? 8'hb1 : _GEN_7509; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7511 = 8'h57 == _t_T_58[7:0] ? 8'h5b : _GEN_7510; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7512 = 8'h58 == _t_T_58[7:0] ? 8'h6a : _GEN_7511; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7513 = 8'h59 == _t_T_58[7:0] ? 8'hcb : _GEN_7512; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7514 = 8'h5a == _t_T_58[7:0] ? 8'hbe : _GEN_7513; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7515 = 8'h5b == _t_T_58[7:0] ? 8'h39 : _GEN_7514; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7516 = 8'h5c == _t_T_58[7:0] ? 8'h4a : _GEN_7515; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7517 = 8'h5d == _t_T_58[7:0] ? 8'h4c : _GEN_7516; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7518 = 8'h5e == _t_T_58[7:0] ? 8'h58 : _GEN_7517; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7519 = 8'h5f == _t_T_58[7:0] ? 8'hcf : _GEN_7518; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7520 = 8'h60 == _t_T_58[7:0] ? 8'hd0 : _GEN_7519; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7521 = 8'h61 == _t_T_58[7:0] ? 8'hef : _GEN_7520; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7522 = 8'h62 == _t_T_58[7:0] ? 8'haa : _GEN_7521; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7523 = 8'h63 == _t_T_58[7:0] ? 8'hfb : _GEN_7522; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7524 = 8'h64 == _t_T_58[7:0] ? 8'h43 : _GEN_7523; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7525 = 8'h65 == _t_T_58[7:0] ? 8'h4d : _GEN_7524; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7526 = 8'h66 == _t_T_58[7:0] ? 8'h33 : _GEN_7525; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7527 = 8'h67 == _t_T_58[7:0] ? 8'h85 : _GEN_7526; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7528 = 8'h68 == _t_T_58[7:0] ? 8'h45 : _GEN_7527; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7529 = 8'h69 == _t_T_58[7:0] ? 8'hf9 : _GEN_7528; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7530 = 8'h6a == _t_T_58[7:0] ? 8'h2 : _GEN_7529; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7531 = 8'h6b == _t_T_58[7:0] ? 8'h7f : _GEN_7530; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7532 = 8'h6c == _t_T_58[7:0] ? 8'h50 : _GEN_7531; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7533 = 8'h6d == _t_T_58[7:0] ? 8'h3c : _GEN_7532; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7534 = 8'h6e == _t_T_58[7:0] ? 8'h9f : _GEN_7533; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7535 = 8'h6f == _t_T_58[7:0] ? 8'ha8 : _GEN_7534; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7536 = 8'h70 == _t_T_58[7:0] ? 8'h51 : _GEN_7535; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7537 = 8'h71 == _t_T_58[7:0] ? 8'ha3 : _GEN_7536; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7538 = 8'h72 == _t_T_58[7:0] ? 8'h40 : _GEN_7537; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7539 = 8'h73 == _t_T_58[7:0] ? 8'h8f : _GEN_7538; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7540 = 8'h74 == _t_T_58[7:0] ? 8'h92 : _GEN_7539; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7541 = 8'h75 == _t_T_58[7:0] ? 8'h9d : _GEN_7540; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7542 = 8'h76 == _t_T_58[7:0] ? 8'h38 : _GEN_7541; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7543 = 8'h77 == _t_T_58[7:0] ? 8'hf5 : _GEN_7542; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7544 = 8'h78 == _t_T_58[7:0] ? 8'hbc : _GEN_7543; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7545 = 8'h79 == _t_T_58[7:0] ? 8'hb6 : _GEN_7544; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7546 = 8'h7a == _t_T_58[7:0] ? 8'hda : _GEN_7545; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7547 = 8'h7b == _t_T_58[7:0] ? 8'h21 : _GEN_7546; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7548 = 8'h7c == _t_T_58[7:0] ? 8'h10 : _GEN_7547; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7549 = 8'h7d == _t_T_58[7:0] ? 8'hff : _GEN_7548; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7550 = 8'h7e == _t_T_58[7:0] ? 8'hf3 : _GEN_7549; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7551 = 8'h7f == _t_T_58[7:0] ? 8'hd2 : _GEN_7550; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7552 = 8'h80 == _t_T_58[7:0] ? 8'hcd : _GEN_7551; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7553 = 8'h81 == _t_T_58[7:0] ? 8'hc : _GEN_7552; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7554 = 8'h82 == _t_T_58[7:0] ? 8'h13 : _GEN_7553; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7555 = 8'h83 == _t_T_58[7:0] ? 8'hec : _GEN_7554; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7556 = 8'h84 == _t_T_58[7:0] ? 8'h5f : _GEN_7555; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7557 = 8'h85 == _t_T_58[7:0] ? 8'h97 : _GEN_7556; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7558 = 8'h86 == _t_T_58[7:0] ? 8'h44 : _GEN_7557; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7559 = 8'h87 == _t_T_58[7:0] ? 8'h17 : _GEN_7558; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7560 = 8'h88 == _t_T_58[7:0] ? 8'hc4 : _GEN_7559; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7561 = 8'h89 == _t_T_58[7:0] ? 8'ha7 : _GEN_7560; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7562 = 8'h8a == _t_T_58[7:0] ? 8'h7e : _GEN_7561; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7563 = 8'h8b == _t_T_58[7:0] ? 8'h3d : _GEN_7562; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7564 = 8'h8c == _t_T_58[7:0] ? 8'h64 : _GEN_7563; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7565 = 8'h8d == _t_T_58[7:0] ? 8'h5d : _GEN_7564; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7566 = 8'h8e == _t_T_58[7:0] ? 8'h19 : _GEN_7565; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7567 = 8'h8f == _t_T_58[7:0] ? 8'h73 : _GEN_7566; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7568 = 8'h90 == _t_T_58[7:0] ? 8'h60 : _GEN_7567; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7569 = 8'h91 == _t_T_58[7:0] ? 8'h81 : _GEN_7568; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7570 = 8'h92 == _t_T_58[7:0] ? 8'h4f : _GEN_7569; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7571 = 8'h93 == _t_T_58[7:0] ? 8'hdc : _GEN_7570; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7572 = 8'h94 == _t_T_58[7:0] ? 8'h22 : _GEN_7571; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7573 = 8'h95 == _t_T_58[7:0] ? 8'h2a : _GEN_7572; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7574 = 8'h96 == _t_T_58[7:0] ? 8'h90 : _GEN_7573; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7575 = 8'h97 == _t_T_58[7:0] ? 8'h88 : _GEN_7574; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7576 = 8'h98 == _t_T_58[7:0] ? 8'h46 : _GEN_7575; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7577 = 8'h99 == _t_T_58[7:0] ? 8'hee : _GEN_7576; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7578 = 8'h9a == _t_T_58[7:0] ? 8'hb8 : _GEN_7577; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7579 = 8'h9b == _t_T_58[7:0] ? 8'h14 : _GEN_7578; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7580 = 8'h9c == _t_T_58[7:0] ? 8'hde : _GEN_7579; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7581 = 8'h9d == _t_T_58[7:0] ? 8'h5e : _GEN_7580; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7582 = 8'h9e == _t_T_58[7:0] ? 8'hb : _GEN_7581; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7583 = 8'h9f == _t_T_58[7:0] ? 8'hdb : _GEN_7582; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7584 = 8'ha0 == _t_T_58[7:0] ? 8'he0 : _GEN_7583; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7585 = 8'ha1 == _t_T_58[7:0] ? 8'h32 : _GEN_7584; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7586 = 8'ha2 == _t_T_58[7:0] ? 8'h3a : _GEN_7585; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7587 = 8'ha3 == _t_T_58[7:0] ? 8'ha : _GEN_7586; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7588 = 8'ha4 == _t_T_58[7:0] ? 8'h49 : _GEN_7587; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7589 = 8'ha5 == _t_T_58[7:0] ? 8'h6 : _GEN_7588; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7590 = 8'ha6 == _t_T_58[7:0] ? 8'h24 : _GEN_7589; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7591 = 8'ha7 == _t_T_58[7:0] ? 8'h5c : _GEN_7590; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7592 = 8'ha8 == _t_T_58[7:0] ? 8'hc2 : _GEN_7591; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7593 = 8'ha9 == _t_T_58[7:0] ? 8'hd3 : _GEN_7592; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7594 = 8'haa == _t_T_58[7:0] ? 8'hac : _GEN_7593; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7595 = 8'hab == _t_T_58[7:0] ? 8'h62 : _GEN_7594; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7596 = 8'hac == _t_T_58[7:0] ? 8'h91 : _GEN_7595; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7597 = 8'had == _t_T_58[7:0] ? 8'h95 : _GEN_7596; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7598 = 8'hae == _t_T_58[7:0] ? 8'he4 : _GEN_7597; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7599 = 8'haf == _t_T_58[7:0] ? 8'h79 : _GEN_7598; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7600 = 8'hb0 == _t_T_58[7:0] ? 8'he7 : _GEN_7599; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7601 = 8'hb1 == _t_T_58[7:0] ? 8'hc8 : _GEN_7600; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7602 = 8'hb2 == _t_T_58[7:0] ? 8'h37 : _GEN_7601; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7603 = 8'hb3 == _t_T_58[7:0] ? 8'h6d : _GEN_7602; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7604 = 8'hb4 == _t_T_58[7:0] ? 8'h8d : _GEN_7603; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7605 = 8'hb5 == _t_T_58[7:0] ? 8'hd5 : _GEN_7604; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7606 = 8'hb6 == _t_T_58[7:0] ? 8'h4e : _GEN_7605; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7607 = 8'hb7 == _t_T_58[7:0] ? 8'ha9 : _GEN_7606; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7608 = 8'hb8 == _t_T_58[7:0] ? 8'h6c : _GEN_7607; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7609 = 8'hb9 == _t_T_58[7:0] ? 8'h56 : _GEN_7608; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7610 = 8'hba == _t_T_58[7:0] ? 8'hf4 : _GEN_7609; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7611 = 8'hbb == _t_T_58[7:0] ? 8'hea : _GEN_7610; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7612 = 8'hbc == _t_T_58[7:0] ? 8'h65 : _GEN_7611; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7613 = 8'hbd == _t_T_58[7:0] ? 8'h7a : _GEN_7612; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7614 = 8'hbe == _t_T_58[7:0] ? 8'hae : _GEN_7613; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7615 = 8'hbf == _t_T_58[7:0] ? 8'h8 : _GEN_7614; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7616 = 8'hc0 == _t_T_58[7:0] ? 8'hba : _GEN_7615; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7617 = 8'hc1 == _t_T_58[7:0] ? 8'h78 : _GEN_7616; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7618 = 8'hc2 == _t_T_58[7:0] ? 8'h25 : _GEN_7617; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7619 = 8'hc3 == _t_T_58[7:0] ? 8'h2e : _GEN_7618; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7620 = 8'hc4 == _t_T_58[7:0] ? 8'h1c : _GEN_7619; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7621 = 8'hc5 == _t_T_58[7:0] ? 8'ha6 : _GEN_7620; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7622 = 8'hc6 == _t_T_58[7:0] ? 8'hb4 : _GEN_7621; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7623 = 8'hc7 == _t_T_58[7:0] ? 8'hc6 : _GEN_7622; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7624 = 8'hc8 == _t_T_58[7:0] ? 8'he8 : _GEN_7623; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7625 = 8'hc9 == _t_T_58[7:0] ? 8'hdd : _GEN_7624; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7626 = 8'hca == _t_T_58[7:0] ? 8'h74 : _GEN_7625; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7627 = 8'hcb == _t_T_58[7:0] ? 8'h1f : _GEN_7626; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7628 = 8'hcc == _t_T_58[7:0] ? 8'h4b : _GEN_7627; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7629 = 8'hcd == _t_T_58[7:0] ? 8'hbd : _GEN_7628; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7630 = 8'hce == _t_T_58[7:0] ? 8'h8b : _GEN_7629; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7631 = 8'hcf == _t_T_58[7:0] ? 8'h8a : _GEN_7630; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7632 = 8'hd0 == _t_T_58[7:0] ? 8'h70 : _GEN_7631; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7633 = 8'hd1 == _t_T_58[7:0] ? 8'h3e : _GEN_7632; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7634 = 8'hd2 == _t_T_58[7:0] ? 8'hb5 : _GEN_7633; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7635 = 8'hd3 == _t_T_58[7:0] ? 8'h66 : _GEN_7634; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7636 = 8'hd4 == _t_T_58[7:0] ? 8'h48 : _GEN_7635; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7637 = 8'hd5 == _t_T_58[7:0] ? 8'h3 : _GEN_7636; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7638 = 8'hd6 == _t_T_58[7:0] ? 8'hf6 : _GEN_7637; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7639 = 8'hd7 == _t_T_58[7:0] ? 8'he : _GEN_7638; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7640 = 8'hd8 == _t_T_58[7:0] ? 8'h61 : _GEN_7639; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7641 = 8'hd9 == _t_T_58[7:0] ? 8'h35 : _GEN_7640; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7642 = 8'hda == _t_T_58[7:0] ? 8'h57 : _GEN_7641; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7643 = 8'hdb == _t_T_58[7:0] ? 8'hb9 : _GEN_7642; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7644 = 8'hdc == _t_T_58[7:0] ? 8'h86 : _GEN_7643; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7645 = 8'hdd == _t_T_58[7:0] ? 8'hc1 : _GEN_7644; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7646 = 8'hde == _t_T_58[7:0] ? 8'h1d : _GEN_7645; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7647 = 8'hdf == _t_T_58[7:0] ? 8'h9e : _GEN_7646; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7648 = 8'he0 == _t_T_58[7:0] ? 8'he1 : _GEN_7647; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7649 = 8'he1 == _t_T_58[7:0] ? 8'hf8 : _GEN_7648; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7650 = 8'he2 == _t_T_58[7:0] ? 8'h98 : _GEN_7649; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7651 = 8'he3 == _t_T_58[7:0] ? 8'h11 : _GEN_7650; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7652 = 8'he4 == _t_T_58[7:0] ? 8'h69 : _GEN_7651; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7653 = 8'he5 == _t_T_58[7:0] ? 8'hd9 : _GEN_7652; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7654 = 8'he6 == _t_T_58[7:0] ? 8'h8e : _GEN_7653; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7655 = 8'he7 == _t_T_58[7:0] ? 8'h94 : _GEN_7654; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7656 = 8'he8 == _t_T_58[7:0] ? 8'h9b : _GEN_7655; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7657 = 8'he9 == _t_T_58[7:0] ? 8'h1e : _GEN_7656; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7658 = 8'hea == _t_T_58[7:0] ? 8'h87 : _GEN_7657; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7659 = 8'heb == _t_T_58[7:0] ? 8'he9 : _GEN_7658; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7660 = 8'hec == _t_T_58[7:0] ? 8'hce : _GEN_7659; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7661 = 8'hed == _t_T_58[7:0] ? 8'h55 : _GEN_7660; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7662 = 8'hee == _t_T_58[7:0] ? 8'h28 : _GEN_7661; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7663 = 8'hef == _t_T_58[7:0] ? 8'hdf : _GEN_7662; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7664 = 8'hf0 == _t_T_58[7:0] ? 8'h8c : _GEN_7663; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7665 = 8'hf1 == _t_T_58[7:0] ? 8'ha1 : _GEN_7664; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7666 = 8'hf2 == _t_T_58[7:0] ? 8'h89 : _GEN_7665; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7667 = 8'hf3 == _t_T_58[7:0] ? 8'hd : _GEN_7666; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7668 = 8'hf4 == _t_T_58[7:0] ? 8'hbf : _GEN_7667; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7669 = 8'hf5 == _t_T_58[7:0] ? 8'he6 : _GEN_7668; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7670 = 8'hf6 == _t_T_58[7:0] ? 8'h42 : _GEN_7669; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7671 = 8'hf7 == _t_T_58[7:0] ? 8'h68 : _GEN_7670; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7672 = 8'hf8 == _t_T_58[7:0] ? 8'h41 : _GEN_7671; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7673 = 8'hf9 == _t_T_58[7:0] ? 8'h99 : _GEN_7672; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7674 = 8'hfa == _t_T_58[7:0] ? 8'h2d : _GEN_7673; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7675 = 8'hfb == _t_T_58[7:0] ? 8'hf : _GEN_7674; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7676 = 8'hfc == _t_T_58[7:0] ? 8'hb0 : _GEN_7675; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7677 = 8'hfd == _t_T_58[7:0] ? 8'h54 : _GEN_7676; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7678 = 8'hfe == _t_T_58[7:0] ? 8'hbb : _GEN_7677; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7679 = 8'hff == _t_T_58[7:0] ? 8'h16 : _GEN_7678; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7681 = 8'h1 == _t_T_58[31:24] ? 8'h7c : 8'h63; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7682 = 8'h2 == _t_T_58[31:24] ? 8'h77 : _GEN_7681; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7683 = 8'h3 == _t_T_58[31:24] ? 8'h7b : _GEN_7682; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7684 = 8'h4 == _t_T_58[31:24] ? 8'hf2 : _GEN_7683; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7685 = 8'h5 == _t_T_58[31:24] ? 8'h6b : _GEN_7684; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7686 = 8'h6 == _t_T_58[31:24] ? 8'h6f : _GEN_7685; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7687 = 8'h7 == _t_T_58[31:24] ? 8'hc5 : _GEN_7686; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7688 = 8'h8 == _t_T_58[31:24] ? 8'h30 : _GEN_7687; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7689 = 8'h9 == _t_T_58[31:24] ? 8'h1 : _GEN_7688; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7690 = 8'ha == _t_T_58[31:24] ? 8'h67 : _GEN_7689; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7691 = 8'hb == _t_T_58[31:24] ? 8'h2b : _GEN_7690; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7692 = 8'hc == _t_T_58[31:24] ? 8'hfe : _GEN_7691; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7693 = 8'hd == _t_T_58[31:24] ? 8'hd7 : _GEN_7692; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7694 = 8'he == _t_T_58[31:24] ? 8'hab : _GEN_7693; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7695 = 8'hf == _t_T_58[31:24] ? 8'h76 : _GEN_7694; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7696 = 8'h10 == _t_T_58[31:24] ? 8'hca : _GEN_7695; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7697 = 8'h11 == _t_T_58[31:24] ? 8'h82 : _GEN_7696; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7698 = 8'h12 == _t_T_58[31:24] ? 8'hc9 : _GEN_7697; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7699 = 8'h13 == _t_T_58[31:24] ? 8'h7d : _GEN_7698; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7700 = 8'h14 == _t_T_58[31:24] ? 8'hfa : _GEN_7699; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7701 = 8'h15 == _t_T_58[31:24] ? 8'h59 : _GEN_7700; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7702 = 8'h16 == _t_T_58[31:24] ? 8'h47 : _GEN_7701; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7703 = 8'h17 == _t_T_58[31:24] ? 8'hf0 : _GEN_7702; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7704 = 8'h18 == _t_T_58[31:24] ? 8'had : _GEN_7703; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7705 = 8'h19 == _t_T_58[31:24] ? 8'hd4 : _GEN_7704; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7706 = 8'h1a == _t_T_58[31:24] ? 8'ha2 : _GEN_7705; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7707 = 8'h1b == _t_T_58[31:24] ? 8'haf : _GEN_7706; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7708 = 8'h1c == _t_T_58[31:24] ? 8'h9c : _GEN_7707; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7709 = 8'h1d == _t_T_58[31:24] ? 8'ha4 : _GEN_7708; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7710 = 8'h1e == _t_T_58[31:24] ? 8'h72 : _GEN_7709; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7711 = 8'h1f == _t_T_58[31:24] ? 8'hc0 : _GEN_7710; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7712 = 8'h20 == _t_T_58[31:24] ? 8'hb7 : _GEN_7711; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7713 = 8'h21 == _t_T_58[31:24] ? 8'hfd : _GEN_7712; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7714 = 8'h22 == _t_T_58[31:24] ? 8'h93 : _GEN_7713; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7715 = 8'h23 == _t_T_58[31:24] ? 8'h26 : _GEN_7714; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7716 = 8'h24 == _t_T_58[31:24] ? 8'h36 : _GEN_7715; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7717 = 8'h25 == _t_T_58[31:24] ? 8'h3f : _GEN_7716; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7718 = 8'h26 == _t_T_58[31:24] ? 8'hf7 : _GEN_7717; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7719 = 8'h27 == _t_T_58[31:24] ? 8'hcc : _GEN_7718; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7720 = 8'h28 == _t_T_58[31:24] ? 8'h34 : _GEN_7719; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7721 = 8'h29 == _t_T_58[31:24] ? 8'ha5 : _GEN_7720; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7722 = 8'h2a == _t_T_58[31:24] ? 8'he5 : _GEN_7721; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7723 = 8'h2b == _t_T_58[31:24] ? 8'hf1 : _GEN_7722; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7724 = 8'h2c == _t_T_58[31:24] ? 8'h71 : _GEN_7723; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7725 = 8'h2d == _t_T_58[31:24] ? 8'hd8 : _GEN_7724; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7726 = 8'h2e == _t_T_58[31:24] ? 8'h31 : _GEN_7725; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7727 = 8'h2f == _t_T_58[31:24] ? 8'h15 : _GEN_7726; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7728 = 8'h30 == _t_T_58[31:24] ? 8'h4 : _GEN_7727; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7729 = 8'h31 == _t_T_58[31:24] ? 8'hc7 : _GEN_7728; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7730 = 8'h32 == _t_T_58[31:24] ? 8'h23 : _GEN_7729; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7731 = 8'h33 == _t_T_58[31:24] ? 8'hc3 : _GEN_7730; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7732 = 8'h34 == _t_T_58[31:24] ? 8'h18 : _GEN_7731; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7733 = 8'h35 == _t_T_58[31:24] ? 8'h96 : _GEN_7732; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7734 = 8'h36 == _t_T_58[31:24] ? 8'h5 : _GEN_7733; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7735 = 8'h37 == _t_T_58[31:24] ? 8'h9a : _GEN_7734; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7736 = 8'h38 == _t_T_58[31:24] ? 8'h7 : _GEN_7735; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7737 = 8'h39 == _t_T_58[31:24] ? 8'h12 : _GEN_7736; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7738 = 8'h3a == _t_T_58[31:24] ? 8'h80 : _GEN_7737; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7739 = 8'h3b == _t_T_58[31:24] ? 8'he2 : _GEN_7738; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7740 = 8'h3c == _t_T_58[31:24] ? 8'heb : _GEN_7739; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7741 = 8'h3d == _t_T_58[31:24] ? 8'h27 : _GEN_7740; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7742 = 8'h3e == _t_T_58[31:24] ? 8'hb2 : _GEN_7741; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7743 = 8'h3f == _t_T_58[31:24] ? 8'h75 : _GEN_7742; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7744 = 8'h40 == _t_T_58[31:24] ? 8'h9 : _GEN_7743; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7745 = 8'h41 == _t_T_58[31:24] ? 8'h83 : _GEN_7744; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7746 = 8'h42 == _t_T_58[31:24] ? 8'h2c : _GEN_7745; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7747 = 8'h43 == _t_T_58[31:24] ? 8'h1a : _GEN_7746; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7748 = 8'h44 == _t_T_58[31:24] ? 8'h1b : _GEN_7747; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7749 = 8'h45 == _t_T_58[31:24] ? 8'h6e : _GEN_7748; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7750 = 8'h46 == _t_T_58[31:24] ? 8'h5a : _GEN_7749; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7751 = 8'h47 == _t_T_58[31:24] ? 8'ha0 : _GEN_7750; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7752 = 8'h48 == _t_T_58[31:24] ? 8'h52 : _GEN_7751; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7753 = 8'h49 == _t_T_58[31:24] ? 8'h3b : _GEN_7752; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7754 = 8'h4a == _t_T_58[31:24] ? 8'hd6 : _GEN_7753; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7755 = 8'h4b == _t_T_58[31:24] ? 8'hb3 : _GEN_7754; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7756 = 8'h4c == _t_T_58[31:24] ? 8'h29 : _GEN_7755; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7757 = 8'h4d == _t_T_58[31:24] ? 8'he3 : _GEN_7756; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7758 = 8'h4e == _t_T_58[31:24] ? 8'h2f : _GEN_7757; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7759 = 8'h4f == _t_T_58[31:24] ? 8'h84 : _GEN_7758; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7760 = 8'h50 == _t_T_58[31:24] ? 8'h53 : _GEN_7759; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7761 = 8'h51 == _t_T_58[31:24] ? 8'hd1 : _GEN_7760; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7762 = 8'h52 == _t_T_58[31:24] ? 8'h0 : _GEN_7761; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7763 = 8'h53 == _t_T_58[31:24] ? 8'hed : _GEN_7762; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7764 = 8'h54 == _t_T_58[31:24] ? 8'h20 : _GEN_7763; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7765 = 8'h55 == _t_T_58[31:24] ? 8'hfc : _GEN_7764; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7766 = 8'h56 == _t_T_58[31:24] ? 8'hb1 : _GEN_7765; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7767 = 8'h57 == _t_T_58[31:24] ? 8'h5b : _GEN_7766; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7768 = 8'h58 == _t_T_58[31:24] ? 8'h6a : _GEN_7767; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7769 = 8'h59 == _t_T_58[31:24] ? 8'hcb : _GEN_7768; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7770 = 8'h5a == _t_T_58[31:24] ? 8'hbe : _GEN_7769; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7771 = 8'h5b == _t_T_58[31:24] ? 8'h39 : _GEN_7770; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7772 = 8'h5c == _t_T_58[31:24] ? 8'h4a : _GEN_7771; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7773 = 8'h5d == _t_T_58[31:24] ? 8'h4c : _GEN_7772; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7774 = 8'h5e == _t_T_58[31:24] ? 8'h58 : _GEN_7773; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7775 = 8'h5f == _t_T_58[31:24] ? 8'hcf : _GEN_7774; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7776 = 8'h60 == _t_T_58[31:24] ? 8'hd0 : _GEN_7775; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7777 = 8'h61 == _t_T_58[31:24] ? 8'hef : _GEN_7776; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7778 = 8'h62 == _t_T_58[31:24] ? 8'haa : _GEN_7777; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7779 = 8'h63 == _t_T_58[31:24] ? 8'hfb : _GEN_7778; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7780 = 8'h64 == _t_T_58[31:24] ? 8'h43 : _GEN_7779; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7781 = 8'h65 == _t_T_58[31:24] ? 8'h4d : _GEN_7780; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7782 = 8'h66 == _t_T_58[31:24] ? 8'h33 : _GEN_7781; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7783 = 8'h67 == _t_T_58[31:24] ? 8'h85 : _GEN_7782; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7784 = 8'h68 == _t_T_58[31:24] ? 8'h45 : _GEN_7783; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7785 = 8'h69 == _t_T_58[31:24] ? 8'hf9 : _GEN_7784; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7786 = 8'h6a == _t_T_58[31:24] ? 8'h2 : _GEN_7785; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7787 = 8'h6b == _t_T_58[31:24] ? 8'h7f : _GEN_7786; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7788 = 8'h6c == _t_T_58[31:24] ? 8'h50 : _GEN_7787; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7789 = 8'h6d == _t_T_58[31:24] ? 8'h3c : _GEN_7788; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7790 = 8'h6e == _t_T_58[31:24] ? 8'h9f : _GEN_7789; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7791 = 8'h6f == _t_T_58[31:24] ? 8'ha8 : _GEN_7790; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7792 = 8'h70 == _t_T_58[31:24] ? 8'h51 : _GEN_7791; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7793 = 8'h71 == _t_T_58[31:24] ? 8'ha3 : _GEN_7792; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7794 = 8'h72 == _t_T_58[31:24] ? 8'h40 : _GEN_7793; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7795 = 8'h73 == _t_T_58[31:24] ? 8'h8f : _GEN_7794; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7796 = 8'h74 == _t_T_58[31:24] ? 8'h92 : _GEN_7795; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7797 = 8'h75 == _t_T_58[31:24] ? 8'h9d : _GEN_7796; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7798 = 8'h76 == _t_T_58[31:24] ? 8'h38 : _GEN_7797; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7799 = 8'h77 == _t_T_58[31:24] ? 8'hf5 : _GEN_7798; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7800 = 8'h78 == _t_T_58[31:24] ? 8'hbc : _GEN_7799; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7801 = 8'h79 == _t_T_58[31:24] ? 8'hb6 : _GEN_7800; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7802 = 8'h7a == _t_T_58[31:24] ? 8'hda : _GEN_7801; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7803 = 8'h7b == _t_T_58[31:24] ? 8'h21 : _GEN_7802; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7804 = 8'h7c == _t_T_58[31:24] ? 8'h10 : _GEN_7803; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7805 = 8'h7d == _t_T_58[31:24] ? 8'hff : _GEN_7804; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7806 = 8'h7e == _t_T_58[31:24] ? 8'hf3 : _GEN_7805; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7807 = 8'h7f == _t_T_58[31:24] ? 8'hd2 : _GEN_7806; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7808 = 8'h80 == _t_T_58[31:24] ? 8'hcd : _GEN_7807; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7809 = 8'h81 == _t_T_58[31:24] ? 8'hc : _GEN_7808; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7810 = 8'h82 == _t_T_58[31:24] ? 8'h13 : _GEN_7809; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7811 = 8'h83 == _t_T_58[31:24] ? 8'hec : _GEN_7810; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7812 = 8'h84 == _t_T_58[31:24] ? 8'h5f : _GEN_7811; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7813 = 8'h85 == _t_T_58[31:24] ? 8'h97 : _GEN_7812; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7814 = 8'h86 == _t_T_58[31:24] ? 8'h44 : _GEN_7813; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7815 = 8'h87 == _t_T_58[31:24] ? 8'h17 : _GEN_7814; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7816 = 8'h88 == _t_T_58[31:24] ? 8'hc4 : _GEN_7815; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7817 = 8'h89 == _t_T_58[31:24] ? 8'ha7 : _GEN_7816; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7818 = 8'h8a == _t_T_58[31:24] ? 8'h7e : _GEN_7817; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7819 = 8'h8b == _t_T_58[31:24] ? 8'h3d : _GEN_7818; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7820 = 8'h8c == _t_T_58[31:24] ? 8'h64 : _GEN_7819; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7821 = 8'h8d == _t_T_58[31:24] ? 8'h5d : _GEN_7820; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7822 = 8'h8e == _t_T_58[31:24] ? 8'h19 : _GEN_7821; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7823 = 8'h8f == _t_T_58[31:24] ? 8'h73 : _GEN_7822; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7824 = 8'h90 == _t_T_58[31:24] ? 8'h60 : _GEN_7823; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7825 = 8'h91 == _t_T_58[31:24] ? 8'h81 : _GEN_7824; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7826 = 8'h92 == _t_T_58[31:24] ? 8'h4f : _GEN_7825; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7827 = 8'h93 == _t_T_58[31:24] ? 8'hdc : _GEN_7826; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7828 = 8'h94 == _t_T_58[31:24] ? 8'h22 : _GEN_7827; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7829 = 8'h95 == _t_T_58[31:24] ? 8'h2a : _GEN_7828; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7830 = 8'h96 == _t_T_58[31:24] ? 8'h90 : _GEN_7829; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7831 = 8'h97 == _t_T_58[31:24] ? 8'h88 : _GEN_7830; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7832 = 8'h98 == _t_T_58[31:24] ? 8'h46 : _GEN_7831; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7833 = 8'h99 == _t_T_58[31:24] ? 8'hee : _GEN_7832; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7834 = 8'h9a == _t_T_58[31:24] ? 8'hb8 : _GEN_7833; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7835 = 8'h9b == _t_T_58[31:24] ? 8'h14 : _GEN_7834; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7836 = 8'h9c == _t_T_58[31:24] ? 8'hde : _GEN_7835; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7837 = 8'h9d == _t_T_58[31:24] ? 8'h5e : _GEN_7836; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7838 = 8'h9e == _t_T_58[31:24] ? 8'hb : _GEN_7837; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7839 = 8'h9f == _t_T_58[31:24] ? 8'hdb : _GEN_7838; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7840 = 8'ha0 == _t_T_58[31:24] ? 8'he0 : _GEN_7839; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7841 = 8'ha1 == _t_T_58[31:24] ? 8'h32 : _GEN_7840; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7842 = 8'ha2 == _t_T_58[31:24] ? 8'h3a : _GEN_7841; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7843 = 8'ha3 == _t_T_58[31:24] ? 8'ha : _GEN_7842; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7844 = 8'ha4 == _t_T_58[31:24] ? 8'h49 : _GEN_7843; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7845 = 8'ha5 == _t_T_58[31:24] ? 8'h6 : _GEN_7844; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7846 = 8'ha6 == _t_T_58[31:24] ? 8'h24 : _GEN_7845; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7847 = 8'ha7 == _t_T_58[31:24] ? 8'h5c : _GEN_7846; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7848 = 8'ha8 == _t_T_58[31:24] ? 8'hc2 : _GEN_7847; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7849 = 8'ha9 == _t_T_58[31:24] ? 8'hd3 : _GEN_7848; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7850 = 8'haa == _t_T_58[31:24] ? 8'hac : _GEN_7849; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7851 = 8'hab == _t_T_58[31:24] ? 8'h62 : _GEN_7850; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7852 = 8'hac == _t_T_58[31:24] ? 8'h91 : _GEN_7851; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7853 = 8'had == _t_T_58[31:24] ? 8'h95 : _GEN_7852; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7854 = 8'hae == _t_T_58[31:24] ? 8'he4 : _GEN_7853; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7855 = 8'haf == _t_T_58[31:24] ? 8'h79 : _GEN_7854; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7856 = 8'hb0 == _t_T_58[31:24] ? 8'he7 : _GEN_7855; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7857 = 8'hb1 == _t_T_58[31:24] ? 8'hc8 : _GEN_7856; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7858 = 8'hb2 == _t_T_58[31:24] ? 8'h37 : _GEN_7857; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7859 = 8'hb3 == _t_T_58[31:24] ? 8'h6d : _GEN_7858; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7860 = 8'hb4 == _t_T_58[31:24] ? 8'h8d : _GEN_7859; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7861 = 8'hb5 == _t_T_58[31:24] ? 8'hd5 : _GEN_7860; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7862 = 8'hb6 == _t_T_58[31:24] ? 8'h4e : _GEN_7861; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7863 = 8'hb7 == _t_T_58[31:24] ? 8'ha9 : _GEN_7862; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7864 = 8'hb8 == _t_T_58[31:24] ? 8'h6c : _GEN_7863; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7865 = 8'hb9 == _t_T_58[31:24] ? 8'h56 : _GEN_7864; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7866 = 8'hba == _t_T_58[31:24] ? 8'hf4 : _GEN_7865; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7867 = 8'hbb == _t_T_58[31:24] ? 8'hea : _GEN_7866; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7868 = 8'hbc == _t_T_58[31:24] ? 8'h65 : _GEN_7867; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7869 = 8'hbd == _t_T_58[31:24] ? 8'h7a : _GEN_7868; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7870 = 8'hbe == _t_T_58[31:24] ? 8'hae : _GEN_7869; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7871 = 8'hbf == _t_T_58[31:24] ? 8'h8 : _GEN_7870; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7872 = 8'hc0 == _t_T_58[31:24] ? 8'hba : _GEN_7871; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7873 = 8'hc1 == _t_T_58[31:24] ? 8'h78 : _GEN_7872; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7874 = 8'hc2 == _t_T_58[31:24] ? 8'h25 : _GEN_7873; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7875 = 8'hc3 == _t_T_58[31:24] ? 8'h2e : _GEN_7874; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7876 = 8'hc4 == _t_T_58[31:24] ? 8'h1c : _GEN_7875; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7877 = 8'hc5 == _t_T_58[31:24] ? 8'ha6 : _GEN_7876; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7878 = 8'hc6 == _t_T_58[31:24] ? 8'hb4 : _GEN_7877; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7879 = 8'hc7 == _t_T_58[31:24] ? 8'hc6 : _GEN_7878; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7880 = 8'hc8 == _t_T_58[31:24] ? 8'he8 : _GEN_7879; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7881 = 8'hc9 == _t_T_58[31:24] ? 8'hdd : _GEN_7880; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7882 = 8'hca == _t_T_58[31:24] ? 8'h74 : _GEN_7881; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7883 = 8'hcb == _t_T_58[31:24] ? 8'h1f : _GEN_7882; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7884 = 8'hcc == _t_T_58[31:24] ? 8'h4b : _GEN_7883; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7885 = 8'hcd == _t_T_58[31:24] ? 8'hbd : _GEN_7884; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7886 = 8'hce == _t_T_58[31:24] ? 8'h8b : _GEN_7885; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7887 = 8'hcf == _t_T_58[31:24] ? 8'h8a : _GEN_7886; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7888 = 8'hd0 == _t_T_58[31:24] ? 8'h70 : _GEN_7887; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7889 = 8'hd1 == _t_T_58[31:24] ? 8'h3e : _GEN_7888; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7890 = 8'hd2 == _t_T_58[31:24] ? 8'hb5 : _GEN_7889; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7891 = 8'hd3 == _t_T_58[31:24] ? 8'h66 : _GEN_7890; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7892 = 8'hd4 == _t_T_58[31:24] ? 8'h48 : _GEN_7891; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7893 = 8'hd5 == _t_T_58[31:24] ? 8'h3 : _GEN_7892; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7894 = 8'hd6 == _t_T_58[31:24] ? 8'hf6 : _GEN_7893; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7895 = 8'hd7 == _t_T_58[31:24] ? 8'he : _GEN_7894; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7896 = 8'hd8 == _t_T_58[31:24] ? 8'h61 : _GEN_7895; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7897 = 8'hd9 == _t_T_58[31:24] ? 8'h35 : _GEN_7896; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7898 = 8'hda == _t_T_58[31:24] ? 8'h57 : _GEN_7897; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7899 = 8'hdb == _t_T_58[31:24] ? 8'hb9 : _GEN_7898; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7900 = 8'hdc == _t_T_58[31:24] ? 8'h86 : _GEN_7899; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7901 = 8'hdd == _t_T_58[31:24] ? 8'hc1 : _GEN_7900; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7902 = 8'hde == _t_T_58[31:24] ? 8'h1d : _GEN_7901; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7903 = 8'hdf == _t_T_58[31:24] ? 8'h9e : _GEN_7902; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7904 = 8'he0 == _t_T_58[31:24] ? 8'he1 : _GEN_7903; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7905 = 8'he1 == _t_T_58[31:24] ? 8'hf8 : _GEN_7904; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7906 = 8'he2 == _t_T_58[31:24] ? 8'h98 : _GEN_7905; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7907 = 8'he3 == _t_T_58[31:24] ? 8'h11 : _GEN_7906; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7908 = 8'he4 == _t_T_58[31:24] ? 8'h69 : _GEN_7907; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7909 = 8'he5 == _t_T_58[31:24] ? 8'hd9 : _GEN_7908; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7910 = 8'he6 == _t_T_58[31:24] ? 8'h8e : _GEN_7909; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7911 = 8'he7 == _t_T_58[31:24] ? 8'h94 : _GEN_7910; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7912 = 8'he8 == _t_T_58[31:24] ? 8'h9b : _GEN_7911; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7913 = 8'he9 == _t_T_58[31:24] ? 8'h1e : _GEN_7912; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7914 = 8'hea == _t_T_58[31:24] ? 8'h87 : _GEN_7913; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7915 = 8'heb == _t_T_58[31:24] ? 8'he9 : _GEN_7914; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7916 = 8'hec == _t_T_58[31:24] ? 8'hce : _GEN_7915; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7917 = 8'hed == _t_T_58[31:24] ? 8'h55 : _GEN_7916; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7918 = 8'hee == _t_T_58[31:24] ? 8'h28 : _GEN_7917; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7919 = 8'hef == _t_T_58[31:24] ? 8'hdf : _GEN_7918; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7920 = 8'hf0 == _t_T_58[31:24] ? 8'h8c : _GEN_7919; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7921 = 8'hf1 == _t_T_58[31:24] ? 8'ha1 : _GEN_7920; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7922 = 8'hf2 == _t_T_58[31:24] ? 8'h89 : _GEN_7921; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7923 = 8'hf3 == _t_T_58[31:24] ? 8'hd : _GEN_7922; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7924 = 8'hf4 == _t_T_58[31:24] ? 8'hbf : _GEN_7923; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7925 = 8'hf5 == _t_T_58[31:24] ? 8'he6 : _GEN_7924; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7926 = 8'hf6 == _t_T_58[31:24] ? 8'h42 : _GEN_7925; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7927 = 8'hf7 == _t_T_58[31:24] ? 8'h68 : _GEN_7926; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7928 = 8'hf8 == _t_T_58[31:24] ? 8'h41 : _GEN_7927; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7929 = 8'hf9 == _t_T_58[31:24] ? 8'h99 : _GEN_7928; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7930 = 8'hfa == _t_T_58[31:24] ? 8'h2d : _GEN_7929; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7931 = 8'hfb == _t_T_58[31:24] ? 8'hf : _GEN_7930; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7932 = 8'hfc == _t_T_58[31:24] ? 8'hb0 : _GEN_7931; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7933 = 8'hfd == _t_T_58[31:24] ? 8'h54 : _GEN_7932; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7934 = 8'hfe == _t_T_58[31:24] ? 8'hbb : _GEN_7933; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7935 = 8'hff == _t_T_58[31:24] ? 8'h16 : _GEN_7934; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7937 = 8'h1 == _t_T_58[23:16] ? 8'h7c : 8'h63; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7938 = 8'h2 == _t_T_58[23:16] ? 8'h77 : _GEN_7937; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7939 = 8'h3 == _t_T_58[23:16] ? 8'h7b : _GEN_7938; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7940 = 8'h4 == _t_T_58[23:16] ? 8'hf2 : _GEN_7939; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7941 = 8'h5 == _t_T_58[23:16] ? 8'h6b : _GEN_7940; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7942 = 8'h6 == _t_T_58[23:16] ? 8'h6f : _GEN_7941; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7943 = 8'h7 == _t_T_58[23:16] ? 8'hc5 : _GEN_7942; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7944 = 8'h8 == _t_T_58[23:16] ? 8'h30 : _GEN_7943; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7945 = 8'h9 == _t_T_58[23:16] ? 8'h1 : _GEN_7944; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7946 = 8'ha == _t_T_58[23:16] ? 8'h67 : _GEN_7945; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7947 = 8'hb == _t_T_58[23:16] ? 8'h2b : _GEN_7946; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7948 = 8'hc == _t_T_58[23:16] ? 8'hfe : _GEN_7947; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7949 = 8'hd == _t_T_58[23:16] ? 8'hd7 : _GEN_7948; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7950 = 8'he == _t_T_58[23:16] ? 8'hab : _GEN_7949; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7951 = 8'hf == _t_T_58[23:16] ? 8'h76 : _GEN_7950; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7952 = 8'h10 == _t_T_58[23:16] ? 8'hca : _GEN_7951; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7953 = 8'h11 == _t_T_58[23:16] ? 8'h82 : _GEN_7952; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7954 = 8'h12 == _t_T_58[23:16] ? 8'hc9 : _GEN_7953; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7955 = 8'h13 == _t_T_58[23:16] ? 8'h7d : _GEN_7954; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7956 = 8'h14 == _t_T_58[23:16] ? 8'hfa : _GEN_7955; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7957 = 8'h15 == _t_T_58[23:16] ? 8'h59 : _GEN_7956; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7958 = 8'h16 == _t_T_58[23:16] ? 8'h47 : _GEN_7957; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7959 = 8'h17 == _t_T_58[23:16] ? 8'hf0 : _GEN_7958; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7960 = 8'h18 == _t_T_58[23:16] ? 8'had : _GEN_7959; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7961 = 8'h19 == _t_T_58[23:16] ? 8'hd4 : _GEN_7960; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7962 = 8'h1a == _t_T_58[23:16] ? 8'ha2 : _GEN_7961; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7963 = 8'h1b == _t_T_58[23:16] ? 8'haf : _GEN_7962; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7964 = 8'h1c == _t_T_58[23:16] ? 8'h9c : _GEN_7963; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7965 = 8'h1d == _t_T_58[23:16] ? 8'ha4 : _GEN_7964; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7966 = 8'h1e == _t_T_58[23:16] ? 8'h72 : _GEN_7965; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7967 = 8'h1f == _t_T_58[23:16] ? 8'hc0 : _GEN_7966; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7968 = 8'h20 == _t_T_58[23:16] ? 8'hb7 : _GEN_7967; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7969 = 8'h21 == _t_T_58[23:16] ? 8'hfd : _GEN_7968; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7970 = 8'h22 == _t_T_58[23:16] ? 8'h93 : _GEN_7969; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7971 = 8'h23 == _t_T_58[23:16] ? 8'h26 : _GEN_7970; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7972 = 8'h24 == _t_T_58[23:16] ? 8'h36 : _GEN_7971; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7973 = 8'h25 == _t_T_58[23:16] ? 8'h3f : _GEN_7972; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7974 = 8'h26 == _t_T_58[23:16] ? 8'hf7 : _GEN_7973; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7975 = 8'h27 == _t_T_58[23:16] ? 8'hcc : _GEN_7974; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7976 = 8'h28 == _t_T_58[23:16] ? 8'h34 : _GEN_7975; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7977 = 8'h29 == _t_T_58[23:16] ? 8'ha5 : _GEN_7976; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7978 = 8'h2a == _t_T_58[23:16] ? 8'he5 : _GEN_7977; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7979 = 8'h2b == _t_T_58[23:16] ? 8'hf1 : _GEN_7978; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7980 = 8'h2c == _t_T_58[23:16] ? 8'h71 : _GEN_7979; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7981 = 8'h2d == _t_T_58[23:16] ? 8'hd8 : _GEN_7980; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7982 = 8'h2e == _t_T_58[23:16] ? 8'h31 : _GEN_7981; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7983 = 8'h2f == _t_T_58[23:16] ? 8'h15 : _GEN_7982; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7984 = 8'h30 == _t_T_58[23:16] ? 8'h4 : _GEN_7983; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7985 = 8'h31 == _t_T_58[23:16] ? 8'hc7 : _GEN_7984; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7986 = 8'h32 == _t_T_58[23:16] ? 8'h23 : _GEN_7985; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7987 = 8'h33 == _t_T_58[23:16] ? 8'hc3 : _GEN_7986; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7988 = 8'h34 == _t_T_58[23:16] ? 8'h18 : _GEN_7987; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7989 = 8'h35 == _t_T_58[23:16] ? 8'h96 : _GEN_7988; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7990 = 8'h36 == _t_T_58[23:16] ? 8'h5 : _GEN_7989; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7991 = 8'h37 == _t_T_58[23:16] ? 8'h9a : _GEN_7990; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7992 = 8'h38 == _t_T_58[23:16] ? 8'h7 : _GEN_7991; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7993 = 8'h39 == _t_T_58[23:16] ? 8'h12 : _GEN_7992; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7994 = 8'h3a == _t_T_58[23:16] ? 8'h80 : _GEN_7993; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7995 = 8'h3b == _t_T_58[23:16] ? 8'he2 : _GEN_7994; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7996 = 8'h3c == _t_T_58[23:16] ? 8'heb : _GEN_7995; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7997 = 8'h3d == _t_T_58[23:16] ? 8'h27 : _GEN_7996; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7998 = 8'h3e == _t_T_58[23:16] ? 8'hb2 : _GEN_7997; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_7999 = 8'h3f == _t_T_58[23:16] ? 8'h75 : _GEN_7998; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8000 = 8'h40 == _t_T_58[23:16] ? 8'h9 : _GEN_7999; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8001 = 8'h41 == _t_T_58[23:16] ? 8'h83 : _GEN_8000; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8002 = 8'h42 == _t_T_58[23:16] ? 8'h2c : _GEN_8001; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8003 = 8'h43 == _t_T_58[23:16] ? 8'h1a : _GEN_8002; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8004 = 8'h44 == _t_T_58[23:16] ? 8'h1b : _GEN_8003; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8005 = 8'h45 == _t_T_58[23:16] ? 8'h6e : _GEN_8004; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8006 = 8'h46 == _t_T_58[23:16] ? 8'h5a : _GEN_8005; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8007 = 8'h47 == _t_T_58[23:16] ? 8'ha0 : _GEN_8006; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8008 = 8'h48 == _t_T_58[23:16] ? 8'h52 : _GEN_8007; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8009 = 8'h49 == _t_T_58[23:16] ? 8'h3b : _GEN_8008; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8010 = 8'h4a == _t_T_58[23:16] ? 8'hd6 : _GEN_8009; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8011 = 8'h4b == _t_T_58[23:16] ? 8'hb3 : _GEN_8010; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8012 = 8'h4c == _t_T_58[23:16] ? 8'h29 : _GEN_8011; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8013 = 8'h4d == _t_T_58[23:16] ? 8'he3 : _GEN_8012; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8014 = 8'h4e == _t_T_58[23:16] ? 8'h2f : _GEN_8013; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8015 = 8'h4f == _t_T_58[23:16] ? 8'h84 : _GEN_8014; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8016 = 8'h50 == _t_T_58[23:16] ? 8'h53 : _GEN_8015; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8017 = 8'h51 == _t_T_58[23:16] ? 8'hd1 : _GEN_8016; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8018 = 8'h52 == _t_T_58[23:16] ? 8'h0 : _GEN_8017; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8019 = 8'h53 == _t_T_58[23:16] ? 8'hed : _GEN_8018; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8020 = 8'h54 == _t_T_58[23:16] ? 8'h20 : _GEN_8019; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8021 = 8'h55 == _t_T_58[23:16] ? 8'hfc : _GEN_8020; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8022 = 8'h56 == _t_T_58[23:16] ? 8'hb1 : _GEN_8021; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8023 = 8'h57 == _t_T_58[23:16] ? 8'h5b : _GEN_8022; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8024 = 8'h58 == _t_T_58[23:16] ? 8'h6a : _GEN_8023; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8025 = 8'h59 == _t_T_58[23:16] ? 8'hcb : _GEN_8024; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8026 = 8'h5a == _t_T_58[23:16] ? 8'hbe : _GEN_8025; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8027 = 8'h5b == _t_T_58[23:16] ? 8'h39 : _GEN_8026; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8028 = 8'h5c == _t_T_58[23:16] ? 8'h4a : _GEN_8027; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8029 = 8'h5d == _t_T_58[23:16] ? 8'h4c : _GEN_8028; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8030 = 8'h5e == _t_T_58[23:16] ? 8'h58 : _GEN_8029; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8031 = 8'h5f == _t_T_58[23:16] ? 8'hcf : _GEN_8030; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8032 = 8'h60 == _t_T_58[23:16] ? 8'hd0 : _GEN_8031; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8033 = 8'h61 == _t_T_58[23:16] ? 8'hef : _GEN_8032; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8034 = 8'h62 == _t_T_58[23:16] ? 8'haa : _GEN_8033; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8035 = 8'h63 == _t_T_58[23:16] ? 8'hfb : _GEN_8034; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8036 = 8'h64 == _t_T_58[23:16] ? 8'h43 : _GEN_8035; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8037 = 8'h65 == _t_T_58[23:16] ? 8'h4d : _GEN_8036; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8038 = 8'h66 == _t_T_58[23:16] ? 8'h33 : _GEN_8037; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8039 = 8'h67 == _t_T_58[23:16] ? 8'h85 : _GEN_8038; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8040 = 8'h68 == _t_T_58[23:16] ? 8'h45 : _GEN_8039; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8041 = 8'h69 == _t_T_58[23:16] ? 8'hf9 : _GEN_8040; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8042 = 8'h6a == _t_T_58[23:16] ? 8'h2 : _GEN_8041; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8043 = 8'h6b == _t_T_58[23:16] ? 8'h7f : _GEN_8042; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8044 = 8'h6c == _t_T_58[23:16] ? 8'h50 : _GEN_8043; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8045 = 8'h6d == _t_T_58[23:16] ? 8'h3c : _GEN_8044; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8046 = 8'h6e == _t_T_58[23:16] ? 8'h9f : _GEN_8045; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8047 = 8'h6f == _t_T_58[23:16] ? 8'ha8 : _GEN_8046; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8048 = 8'h70 == _t_T_58[23:16] ? 8'h51 : _GEN_8047; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8049 = 8'h71 == _t_T_58[23:16] ? 8'ha3 : _GEN_8048; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8050 = 8'h72 == _t_T_58[23:16] ? 8'h40 : _GEN_8049; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8051 = 8'h73 == _t_T_58[23:16] ? 8'h8f : _GEN_8050; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8052 = 8'h74 == _t_T_58[23:16] ? 8'h92 : _GEN_8051; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8053 = 8'h75 == _t_T_58[23:16] ? 8'h9d : _GEN_8052; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8054 = 8'h76 == _t_T_58[23:16] ? 8'h38 : _GEN_8053; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8055 = 8'h77 == _t_T_58[23:16] ? 8'hf5 : _GEN_8054; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8056 = 8'h78 == _t_T_58[23:16] ? 8'hbc : _GEN_8055; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8057 = 8'h79 == _t_T_58[23:16] ? 8'hb6 : _GEN_8056; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8058 = 8'h7a == _t_T_58[23:16] ? 8'hda : _GEN_8057; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8059 = 8'h7b == _t_T_58[23:16] ? 8'h21 : _GEN_8058; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8060 = 8'h7c == _t_T_58[23:16] ? 8'h10 : _GEN_8059; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8061 = 8'h7d == _t_T_58[23:16] ? 8'hff : _GEN_8060; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8062 = 8'h7e == _t_T_58[23:16] ? 8'hf3 : _GEN_8061; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8063 = 8'h7f == _t_T_58[23:16] ? 8'hd2 : _GEN_8062; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8064 = 8'h80 == _t_T_58[23:16] ? 8'hcd : _GEN_8063; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8065 = 8'h81 == _t_T_58[23:16] ? 8'hc : _GEN_8064; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8066 = 8'h82 == _t_T_58[23:16] ? 8'h13 : _GEN_8065; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8067 = 8'h83 == _t_T_58[23:16] ? 8'hec : _GEN_8066; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8068 = 8'h84 == _t_T_58[23:16] ? 8'h5f : _GEN_8067; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8069 = 8'h85 == _t_T_58[23:16] ? 8'h97 : _GEN_8068; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8070 = 8'h86 == _t_T_58[23:16] ? 8'h44 : _GEN_8069; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8071 = 8'h87 == _t_T_58[23:16] ? 8'h17 : _GEN_8070; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8072 = 8'h88 == _t_T_58[23:16] ? 8'hc4 : _GEN_8071; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8073 = 8'h89 == _t_T_58[23:16] ? 8'ha7 : _GEN_8072; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8074 = 8'h8a == _t_T_58[23:16] ? 8'h7e : _GEN_8073; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8075 = 8'h8b == _t_T_58[23:16] ? 8'h3d : _GEN_8074; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8076 = 8'h8c == _t_T_58[23:16] ? 8'h64 : _GEN_8075; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8077 = 8'h8d == _t_T_58[23:16] ? 8'h5d : _GEN_8076; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8078 = 8'h8e == _t_T_58[23:16] ? 8'h19 : _GEN_8077; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8079 = 8'h8f == _t_T_58[23:16] ? 8'h73 : _GEN_8078; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8080 = 8'h90 == _t_T_58[23:16] ? 8'h60 : _GEN_8079; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8081 = 8'h91 == _t_T_58[23:16] ? 8'h81 : _GEN_8080; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8082 = 8'h92 == _t_T_58[23:16] ? 8'h4f : _GEN_8081; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8083 = 8'h93 == _t_T_58[23:16] ? 8'hdc : _GEN_8082; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8084 = 8'h94 == _t_T_58[23:16] ? 8'h22 : _GEN_8083; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8085 = 8'h95 == _t_T_58[23:16] ? 8'h2a : _GEN_8084; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8086 = 8'h96 == _t_T_58[23:16] ? 8'h90 : _GEN_8085; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8087 = 8'h97 == _t_T_58[23:16] ? 8'h88 : _GEN_8086; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8088 = 8'h98 == _t_T_58[23:16] ? 8'h46 : _GEN_8087; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8089 = 8'h99 == _t_T_58[23:16] ? 8'hee : _GEN_8088; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8090 = 8'h9a == _t_T_58[23:16] ? 8'hb8 : _GEN_8089; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8091 = 8'h9b == _t_T_58[23:16] ? 8'h14 : _GEN_8090; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8092 = 8'h9c == _t_T_58[23:16] ? 8'hde : _GEN_8091; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8093 = 8'h9d == _t_T_58[23:16] ? 8'h5e : _GEN_8092; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8094 = 8'h9e == _t_T_58[23:16] ? 8'hb : _GEN_8093; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8095 = 8'h9f == _t_T_58[23:16] ? 8'hdb : _GEN_8094; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8096 = 8'ha0 == _t_T_58[23:16] ? 8'he0 : _GEN_8095; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8097 = 8'ha1 == _t_T_58[23:16] ? 8'h32 : _GEN_8096; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8098 = 8'ha2 == _t_T_58[23:16] ? 8'h3a : _GEN_8097; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8099 = 8'ha3 == _t_T_58[23:16] ? 8'ha : _GEN_8098; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8100 = 8'ha4 == _t_T_58[23:16] ? 8'h49 : _GEN_8099; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8101 = 8'ha5 == _t_T_58[23:16] ? 8'h6 : _GEN_8100; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8102 = 8'ha6 == _t_T_58[23:16] ? 8'h24 : _GEN_8101; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8103 = 8'ha7 == _t_T_58[23:16] ? 8'h5c : _GEN_8102; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8104 = 8'ha8 == _t_T_58[23:16] ? 8'hc2 : _GEN_8103; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8105 = 8'ha9 == _t_T_58[23:16] ? 8'hd3 : _GEN_8104; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8106 = 8'haa == _t_T_58[23:16] ? 8'hac : _GEN_8105; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8107 = 8'hab == _t_T_58[23:16] ? 8'h62 : _GEN_8106; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8108 = 8'hac == _t_T_58[23:16] ? 8'h91 : _GEN_8107; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8109 = 8'had == _t_T_58[23:16] ? 8'h95 : _GEN_8108; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8110 = 8'hae == _t_T_58[23:16] ? 8'he4 : _GEN_8109; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8111 = 8'haf == _t_T_58[23:16] ? 8'h79 : _GEN_8110; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8112 = 8'hb0 == _t_T_58[23:16] ? 8'he7 : _GEN_8111; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8113 = 8'hb1 == _t_T_58[23:16] ? 8'hc8 : _GEN_8112; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8114 = 8'hb2 == _t_T_58[23:16] ? 8'h37 : _GEN_8113; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8115 = 8'hb3 == _t_T_58[23:16] ? 8'h6d : _GEN_8114; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8116 = 8'hb4 == _t_T_58[23:16] ? 8'h8d : _GEN_8115; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8117 = 8'hb5 == _t_T_58[23:16] ? 8'hd5 : _GEN_8116; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8118 = 8'hb6 == _t_T_58[23:16] ? 8'h4e : _GEN_8117; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8119 = 8'hb7 == _t_T_58[23:16] ? 8'ha9 : _GEN_8118; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8120 = 8'hb8 == _t_T_58[23:16] ? 8'h6c : _GEN_8119; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8121 = 8'hb9 == _t_T_58[23:16] ? 8'h56 : _GEN_8120; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8122 = 8'hba == _t_T_58[23:16] ? 8'hf4 : _GEN_8121; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8123 = 8'hbb == _t_T_58[23:16] ? 8'hea : _GEN_8122; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8124 = 8'hbc == _t_T_58[23:16] ? 8'h65 : _GEN_8123; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8125 = 8'hbd == _t_T_58[23:16] ? 8'h7a : _GEN_8124; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8126 = 8'hbe == _t_T_58[23:16] ? 8'hae : _GEN_8125; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8127 = 8'hbf == _t_T_58[23:16] ? 8'h8 : _GEN_8126; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8128 = 8'hc0 == _t_T_58[23:16] ? 8'hba : _GEN_8127; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8129 = 8'hc1 == _t_T_58[23:16] ? 8'h78 : _GEN_8128; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8130 = 8'hc2 == _t_T_58[23:16] ? 8'h25 : _GEN_8129; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8131 = 8'hc3 == _t_T_58[23:16] ? 8'h2e : _GEN_8130; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8132 = 8'hc4 == _t_T_58[23:16] ? 8'h1c : _GEN_8131; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8133 = 8'hc5 == _t_T_58[23:16] ? 8'ha6 : _GEN_8132; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8134 = 8'hc6 == _t_T_58[23:16] ? 8'hb4 : _GEN_8133; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8135 = 8'hc7 == _t_T_58[23:16] ? 8'hc6 : _GEN_8134; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8136 = 8'hc8 == _t_T_58[23:16] ? 8'he8 : _GEN_8135; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8137 = 8'hc9 == _t_T_58[23:16] ? 8'hdd : _GEN_8136; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8138 = 8'hca == _t_T_58[23:16] ? 8'h74 : _GEN_8137; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8139 = 8'hcb == _t_T_58[23:16] ? 8'h1f : _GEN_8138; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8140 = 8'hcc == _t_T_58[23:16] ? 8'h4b : _GEN_8139; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8141 = 8'hcd == _t_T_58[23:16] ? 8'hbd : _GEN_8140; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8142 = 8'hce == _t_T_58[23:16] ? 8'h8b : _GEN_8141; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8143 = 8'hcf == _t_T_58[23:16] ? 8'h8a : _GEN_8142; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8144 = 8'hd0 == _t_T_58[23:16] ? 8'h70 : _GEN_8143; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8145 = 8'hd1 == _t_T_58[23:16] ? 8'h3e : _GEN_8144; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8146 = 8'hd2 == _t_T_58[23:16] ? 8'hb5 : _GEN_8145; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8147 = 8'hd3 == _t_T_58[23:16] ? 8'h66 : _GEN_8146; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8148 = 8'hd4 == _t_T_58[23:16] ? 8'h48 : _GEN_8147; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8149 = 8'hd5 == _t_T_58[23:16] ? 8'h3 : _GEN_8148; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8150 = 8'hd6 == _t_T_58[23:16] ? 8'hf6 : _GEN_8149; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8151 = 8'hd7 == _t_T_58[23:16] ? 8'he : _GEN_8150; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8152 = 8'hd8 == _t_T_58[23:16] ? 8'h61 : _GEN_8151; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8153 = 8'hd9 == _t_T_58[23:16] ? 8'h35 : _GEN_8152; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8154 = 8'hda == _t_T_58[23:16] ? 8'h57 : _GEN_8153; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8155 = 8'hdb == _t_T_58[23:16] ? 8'hb9 : _GEN_8154; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8156 = 8'hdc == _t_T_58[23:16] ? 8'h86 : _GEN_8155; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8157 = 8'hdd == _t_T_58[23:16] ? 8'hc1 : _GEN_8156; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8158 = 8'hde == _t_T_58[23:16] ? 8'h1d : _GEN_8157; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8159 = 8'hdf == _t_T_58[23:16] ? 8'h9e : _GEN_8158; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8160 = 8'he0 == _t_T_58[23:16] ? 8'he1 : _GEN_8159; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8161 = 8'he1 == _t_T_58[23:16] ? 8'hf8 : _GEN_8160; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8162 = 8'he2 == _t_T_58[23:16] ? 8'h98 : _GEN_8161; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8163 = 8'he3 == _t_T_58[23:16] ? 8'h11 : _GEN_8162; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8164 = 8'he4 == _t_T_58[23:16] ? 8'h69 : _GEN_8163; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8165 = 8'he5 == _t_T_58[23:16] ? 8'hd9 : _GEN_8164; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8166 = 8'he6 == _t_T_58[23:16] ? 8'h8e : _GEN_8165; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8167 = 8'he7 == _t_T_58[23:16] ? 8'h94 : _GEN_8166; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8168 = 8'he8 == _t_T_58[23:16] ? 8'h9b : _GEN_8167; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8169 = 8'he9 == _t_T_58[23:16] ? 8'h1e : _GEN_8168; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8170 = 8'hea == _t_T_58[23:16] ? 8'h87 : _GEN_8169; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8171 = 8'heb == _t_T_58[23:16] ? 8'he9 : _GEN_8170; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8172 = 8'hec == _t_T_58[23:16] ? 8'hce : _GEN_8171; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8173 = 8'hed == _t_T_58[23:16] ? 8'h55 : _GEN_8172; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8174 = 8'hee == _t_T_58[23:16] ? 8'h28 : _GEN_8173; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8175 = 8'hef == _t_T_58[23:16] ? 8'hdf : _GEN_8174; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8176 = 8'hf0 == _t_T_58[23:16] ? 8'h8c : _GEN_8175; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8177 = 8'hf1 == _t_T_58[23:16] ? 8'ha1 : _GEN_8176; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8178 = 8'hf2 == _t_T_58[23:16] ? 8'h89 : _GEN_8177; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8179 = 8'hf3 == _t_T_58[23:16] ? 8'hd : _GEN_8178; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8180 = 8'hf4 == _t_T_58[23:16] ? 8'hbf : _GEN_8179; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8181 = 8'hf5 == _t_T_58[23:16] ? 8'he6 : _GEN_8180; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8182 = 8'hf6 == _t_T_58[23:16] ? 8'h42 : _GEN_8181; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8183 = 8'hf7 == _t_T_58[23:16] ? 8'h68 : _GEN_8182; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8184 = 8'hf8 == _t_T_58[23:16] ? 8'h41 : _GEN_8183; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8185 = 8'hf9 == _t_T_58[23:16] ? 8'h99 : _GEN_8184; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8186 = 8'hfa == _t_T_58[23:16] ? 8'h2d : _GEN_8185; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8187 = 8'hfb == _t_T_58[23:16] ? 8'hf : _GEN_8186; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8188 = 8'hfc == _t_T_58[23:16] ? 8'hb0 : _GEN_8187; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8189 = 8'hfd == _t_T_58[23:16] ? 8'h54 : _GEN_8188; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8190 = 8'hfe == _t_T_58[23:16] ? 8'hbb : _GEN_8189; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8191 = 8'hff == _t_T_58[23:16] ? 8'h16 : _GEN_8190; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [31:0] _t_T_63 = {_GEN_7935,_GEN_8191,_GEN_7423,_GEN_7679}; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:8]
  wire [31:0] t_7 = _t_T_63 ^ 32'h80000000; // @[src/main/scala/crypto/aes/KeySchedule.scala 59:32]
  wire [31:0] w_32 = w_28 ^ t_7; // @[src/main/scala/crypto/aes/KeySchedule.scala 63:21]
  wire [31:0] w_33 = w_29 ^ w_32; // @[src/main/scala/crypto/aes/KeySchedule.scala 63:21]
  wire [31:0] w_34 = w_30 ^ w_33; // @[src/main/scala/crypto/aes/KeySchedule.scala 63:21]
  wire [31:0] w_35 = w_31 ^ w_34; // @[src/main/scala/crypto/aes/KeySchedule.scala 63:21]
  wire [31:0] _t_T_66 = {w_35[23:0],w_35[31:24]}; // @[src/main/scala/crypto/aes/KeySchedule.scala 23:43]
  wire [7:0] _GEN_8193 = 8'h1 == _t_T_66[15:8] ? 8'h7c : 8'h63; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8194 = 8'h2 == _t_T_66[15:8] ? 8'h77 : _GEN_8193; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8195 = 8'h3 == _t_T_66[15:8] ? 8'h7b : _GEN_8194; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8196 = 8'h4 == _t_T_66[15:8] ? 8'hf2 : _GEN_8195; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8197 = 8'h5 == _t_T_66[15:8] ? 8'h6b : _GEN_8196; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8198 = 8'h6 == _t_T_66[15:8] ? 8'h6f : _GEN_8197; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8199 = 8'h7 == _t_T_66[15:8] ? 8'hc5 : _GEN_8198; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8200 = 8'h8 == _t_T_66[15:8] ? 8'h30 : _GEN_8199; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8201 = 8'h9 == _t_T_66[15:8] ? 8'h1 : _GEN_8200; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8202 = 8'ha == _t_T_66[15:8] ? 8'h67 : _GEN_8201; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8203 = 8'hb == _t_T_66[15:8] ? 8'h2b : _GEN_8202; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8204 = 8'hc == _t_T_66[15:8] ? 8'hfe : _GEN_8203; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8205 = 8'hd == _t_T_66[15:8] ? 8'hd7 : _GEN_8204; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8206 = 8'he == _t_T_66[15:8] ? 8'hab : _GEN_8205; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8207 = 8'hf == _t_T_66[15:8] ? 8'h76 : _GEN_8206; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8208 = 8'h10 == _t_T_66[15:8] ? 8'hca : _GEN_8207; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8209 = 8'h11 == _t_T_66[15:8] ? 8'h82 : _GEN_8208; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8210 = 8'h12 == _t_T_66[15:8] ? 8'hc9 : _GEN_8209; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8211 = 8'h13 == _t_T_66[15:8] ? 8'h7d : _GEN_8210; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8212 = 8'h14 == _t_T_66[15:8] ? 8'hfa : _GEN_8211; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8213 = 8'h15 == _t_T_66[15:8] ? 8'h59 : _GEN_8212; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8214 = 8'h16 == _t_T_66[15:8] ? 8'h47 : _GEN_8213; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8215 = 8'h17 == _t_T_66[15:8] ? 8'hf0 : _GEN_8214; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8216 = 8'h18 == _t_T_66[15:8] ? 8'had : _GEN_8215; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8217 = 8'h19 == _t_T_66[15:8] ? 8'hd4 : _GEN_8216; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8218 = 8'h1a == _t_T_66[15:8] ? 8'ha2 : _GEN_8217; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8219 = 8'h1b == _t_T_66[15:8] ? 8'haf : _GEN_8218; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8220 = 8'h1c == _t_T_66[15:8] ? 8'h9c : _GEN_8219; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8221 = 8'h1d == _t_T_66[15:8] ? 8'ha4 : _GEN_8220; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8222 = 8'h1e == _t_T_66[15:8] ? 8'h72 : _GEN_8221; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8223 = 8'h1f == _t_T_66[15:8] ? 8'hc0 : _GEN_8222; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8224 = 8'h20 == _t_T_66[15:8] ? 8'hb7 : _GEN_8223; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8225 = 8'h21 == _t_T_66[15:8] ? 8'hfd : _GEN_8224; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8226 = 8'h22 == _t_T_66[15:8] ? 8'h93 : _GEN_8225; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8227 = 8'h23 == _t_T_66[15:8] ? 8'h26 : _GEN_8226; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8228 = 8'h24 == _t_T_66[15:8] ? 8'h36 : _GEN_8227; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8229 = 8'h25 == _t_T_66[15:8] ? 8'h3f : _GEN_8228; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8230 = 8'h26 == _t_T_66[15:8] ? 8'hf7 : _GEN_8229; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8231 = 8'h27 == _t_T_66[15:8] ? 8'hcc : _GEN_8230; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8232 = 8'h28 == _t_T_66[15:8] ? 8'h34 : _GEN_8231; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8233 = 8'h29 == _t_T_66[15:8] ? 8'ha5 : _GEN_8232; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8234 = 8'h2a == _t_T_66[15:8] ? 8'he5 : _GEN_8233; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8235 = 8'h2b == _t_T_66[15:8] ? 8'hf1 : _GEN_8234; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8236 = 8'h2c == _t_T_66[15:8] ? 8'h71 : _GEN_8235; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8237 = 8'h2d == _t_T_66[15:8] ? 8'hd8 : _GEN_8236; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8238 = 8'h2e == _t_T_66[15:8] ? 8'h31 : _GEN_8237; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8239 = 8'h2f == _t_T_66[15:8] ? 8'h15 : _GEN_8238; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8240 = 8'h30 == _t_T_66[15:8] ? 8'h4 : _GEN_8239; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8241 = 8'h31 == _t_T_66[15:8] ? 8'hc7 : _GEN_8240; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8242 = 8'h32 == _t_T_66[15:8] ? 8'h23 : _GEN_8241; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8243 = 8'h33 == _t_T_66[15:8] ? 8'hc3 : _GEN_8242; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8244 = 8'h34 == _t_T_66[15:8] ? 8'h18 : _GEN_8243; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8245 = 8'h35 == _t_T_66[15:8] ? 8'h96 : _GEN_8244; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8246 = 8'h36 == _t_T_66[15:8] ? 8'h5 : _GEN_8245; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8247 = 8'h37 == _t_T_66[15:8] ? 8'h9a : _GEN_8246; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8248 = 8'h38 == _t_T_66[15:8] ? 8'h7 : _GEN_8247; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8249 = 8'h39 == _t_T_66[15:8] ? 8'h12 : _GEN_8248; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8250 = 8'h3a == _t_T_66[15:8] ? 8'h80 : _GEN_8249; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8251 = 8'h3b == _t_T_66[15:8] ? 8'he2 : _GEN_8250; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8252 = 8'h3c == _t_T_66[15:8] ? 8'heb : _GEN_8251; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8253 = 8'h3d == _t_T_66[15:8] ? 8'h27 : _GEN_8252; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8254 = 8'h3e == _t_T_66[15:8] ? 8'hb2 : _GEN_8253; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8255 = 8'h3f == _t_T_66[15:8] ? 8'h75 : _GEN_8254; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8256 = 8'h40 == _t_T_66[15:8] ? 8'h9 : _GEN_8255; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8257 = 8'h41 == _t_T_66[15:8] ? 8'h83 : _GEN_8256; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8258 = 8'h42 == _t_T_66[15:8] ? 8'h2c : _GEN_8257; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8259 = 8'h43 == _t_T_66[15:8] ? 8'h1a : _GEN_8258; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8260 = 8'h44 == _t_T_66[15:8] ? 8'h1b : _GEN_8259; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8261 = 8'h45 == _t_T_66[15:8] ? 8'h6e : _GEN_8260; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8262 = 8'h46 == _t_T_66[15:8] ? 8'h5a : _GEN_8261; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8263 = 8'h47 == _t_T_66[15:8] ? 8'ha0 : _GEN_8262; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8264 = 8'h48 == _t_T_66[15:8] ? 8'h52 : _GEN_8263; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8265 = 8'h49 == _t_T_66[15:8] ? 8'h3b : _GEN_8264; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8266 = 8'h4a == _t_T_66[15:8] ? 8'hd6 : _GEN_8265; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8267 = 8'h4b == _t_T_66[15:8] ? 8'hb3 : _GEN_8266; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8268 = 8'h4c == _t_T_66[15:8] ? 8'h29 : _GEN_8267; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8269 = 8'h4d == _t_T_66[15:8] ? 8'he3 : _GEN_8268; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8270 = 8'h4e == _t_T_66[15:8] ? 8'h2f : _GEN_8269; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8271 = 8'h4f == _t_T_66[15:8] ? 8'h84 : _GEN_8270; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8272 = 8'h50 == _t_T_66[15:8] ? 8'h53 : _GEN_8271; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8273 = 8'h51 == _t_T_66[15:8] ? 8'hd1 : _GEN_8272; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8274 = 8'h52 == _t_T_66[15:8] ? 8'h0 : _GEN_8273; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8275 = 8'h53 == _t_T_66[15:8] ? 8'hed : _GEN_8274; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8276 = 8'h54 == _t_T_66[15:8] ? 8'h20 : _GEN_8275; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8277 = 8'h55 == _t_T_66[15:8] ? 8'hfc : _GEN_8276; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8278 = 8'h56 == _t_T_66[15:8] ? 8'hb1 : _GEN_8277; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8279 = 8'h57 == _t_T_66[15:8] ? 8'h5b : _GEN_8278; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8280 = 8'h58 == _t_T_66[15:8] ? 8'h6a : _GEN_8279; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8281 = 8'h59 == _t_T_66[15:8] ? 8'hcb : _GEN_8280; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8282 = 8'h5a == _t_T_66[15:8] ? 8'hbe : _GEN_8281; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8283 = 8'h5b == _t_T_66[15:8] ? 8'h39 : _GEN_8282; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8284 = 8'h5c == _t_T_66[15:8] ? 8'h4a : _GEN_8283; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8285 = 8'h5d == _t_T_66[15:8] ? 8'h4c : _GEN_8284; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8286 = 8'h5e == _t_T_66[15:8] ? 8'h58 : _GEN_8285; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8287 = 8'h5f == _t_T_66[15:8] ? 8'hcf : _GEN_8286; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8288 = 8'h60 == _t_T_66[15:8] ? 8'hd0 : _GEN_8287; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8289 = 8'h61 == _t_T_66[15:8] ? 8'hef : _GEN_8288; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8290 = 8'h62 == _t_T_66[15:8] ? 8'haa : _GEN_8289; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8291 = 8'h63 == _t_T_66[15:8] ? 8'hfb : _GEN_8290; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8292 = 8'h64 == _t_T_66[15:8] ? 8'h43 : _GEN_8291; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8293 = 8'h65 == _t_T_66[15:8] ? 8'h4d : _GEN_8292; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8294 = 8'h66 == _t_T_66[15:8] ? 8'h33 : _GEN_8293; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8295 = 8'h67 == _t_T_66[15:8] ? 8'h85 : _GEN_8294; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8296 = 8'h68 == _t_T_66[15:8] ? 8'h45 : _GEN_8295; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8297 = 8'h69 == _t_T_66[15:8] ? 8'hf9 : _GEN_8296; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8298 = 8'h6a == _t_T_66[15:8] ? 8'h2 : _GEN_8297; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8299 = 8'h6b == _t_T_66[15:8] ? 8'h7f : _GEN_8298; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8300 = 8'h6c == _t_T_66[15:8] ? 8'h50 : _GEN_8299; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8301 = 8'h6d == _t_T_66[15:8] ? 8'h3c : _GEN_8300; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8302 = 8'h6e == _t_T_66[15:8] ? 8'h9f : _GEN_8301; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8303 = 8'h6f == _t_T_66[15:8] ? 8'ha8 : _GEN_8302; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8304 = 8'h70 == _t_T_66[15:8] ? 8'h51 : _GEN_8303; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8305 = 8'h71 == _t_T_66[15:8] ? 8'ha3 : _GEN_8304; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8306 = 8'h72 == _t_T_66[15:8] ? 8'h40 : _GEN_8305; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8307 = 8'h73 == _t_T_66[15:8] ? 8'h8f : _GEN_8306; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8308 = 8'h74 == _t_T_66[15:8] ? 8'h92 : _GEN_8307; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8309 = 8'h75 == _t_T_66[15:8] ? 8'h9d : _GEN_8308; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8310 = 8'h76 == _t_T_66[15:8] ? 8'h38 : _GEN_8309; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8311 = 8'h77 == _t_T_66[15:8] ? 8'hf5 : _GEN_8310; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8312 = 8'h78 == _t_T_66[15:8] ? 8'hbc : _GEN_8311; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8313 = 8'h79 == _t_T_66[15:8] ? 8'hb6 : _GEN_8312; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8314 = 8'h7a == _t_T_66[15:8] ? 8'hda : _GEN_8313; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8315 = 8'h7b == _t_T_66[15:8] ? 8'h21 : _GEN_8314; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8316 = 8'h7c == _t_T_66[15:8] ? 8'h10 : _GEN_8315; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8317 = 8'h7d == _t_T_66[15:8] ? 8'hff : _GEN_8316; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8318 = 8'h7e == _t_T_66[15:8] ? 8'hf3 : _GEN_8317; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8319 = 8'h7f == _t_T_66[15:8] ? 8'hd2 : _GEN_8318; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8320 = 8'h80 == _t_T_66[15:8] ? 8'hcd : _GEN_8319; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8321 = 8'h81 == _t_T_66[15:8] ? 8'hc : _GEN_8320; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8322 = 8'h82 == _t_T_66[15:8] ? 8'h13 : _GEN_8321; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8323 = 8'h83 == _t_T_66[15:8] ? 8'hec : _GEN_8322; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8324 = 8'h84 == _t_T_66[15:8] ? 8'h5f : _GEN_8323; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8325 = 8'h85 == _t_T_66[15:8] ? 8'h97 : _GEN_8324; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8326 = 8'h86 == _t_T_66[15:8] ? 8'h44 : _GEN_8325; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8327 = 8'h87 == _t_T_66[15:8] ? 8'h17 : _GEN_8326; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8328 = 8'h88 == _t_T_66[15:8] ? 8'hc4 : _GEN_8327; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8329 = 8'h89 == _t_T_66[15:8] ? 8'ha7 : _GEN_8328; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8330 = 8'h8a == _t_T_66[15:8] ? 8'h7e : _GEN_8329; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8331 = 8'h8b == _t_T_66[15:8] ? 8'h3d : _GEN_8330; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8332 = 8'h8c == _t_T_66[15:8] ? 8'h64 : _GEN_8331; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8333 = 8'h8d == _t_T_66[15:8] ? 8'h5d : _GEN_8332; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8334 = 8'h8e == _t_T_66[15:8] ? 8'h19 : _GEN_8333; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8335 = 8'h8f == _t_T_66[15:8] ? 8'h73 : _GEN_8334; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8336 = 8'h90 == _t_T_66[15:8] ? 8'h60 : _GEN_8335; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8337 = 8'h91 == _t_T_66[15:8] ? 8'h81 : _GEN_8336; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8338 = 8'h92 == _t_T_66[15:8] ? 8'h4f : _GEN_8337; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8339 = 8'h93 == _t_T_66[15:8] ? 8'hdc : _GEN_8338; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8340 = 8'h94 == _t_T_66[15:8] ? 8'h22 : _GEN_8339; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8341 = 8'h95 == _t_T_66[15:8] ? 8'h2a : _GEN_8340; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8342 = 8'h96 == _t_T_66[15:8] ? 8'h90 : _GEN_8341; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8343 = 8'h97 == _t_T_66[15:8] ? 8'h88 : _GEN_8342; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8344 = 8'h98 == _t_T_66[15:8] ? 8'h46 : _GEN_8343; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8345 = 8'h99 == _t_T_66[15:8] ? 8'hee : _GEN_8344; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8346 = 8'h9a == _t_T_66[15:8] ? 8'hb8 : _GEN_8345; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8347 = 8'h9b == _t_T_66[15:8] ? 8'h14 : _GEN_8346; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8348 = 8'h9c == _t_T_66[15:8] ? 8'hde : _GEN_8347; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8349 = 8'h9d == _t_T_66[15:8] ? 8'h5e : _GEN_8348; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8350 = 8'h9e == _t_T_66[15:8] ? 8'hb : _GEN_8349; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8351 = 8'h9f == _t_T_66[15:8] ? 8'hdb : _GEN_8350; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8352 = 8'ha0 == _t_T_66[15:8] ? 8'he0 : _GEN_8351; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8353 = 8'ha1 == _t_T_66[15:8] ? 8'h32 : _GEN_8352; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8354 = 8'ha2 == _t_T_66[15:8] ? 8'h3a : _GEN_8353; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8355 = 8'ha3 == _t_T_66[15:8] ? 8'ha : _GEN_8354; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8356 = 8'ha4 == _t_T_66[15:8] ? 8'h49 : _GEN_8355; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8357 = 8'ha5 == _t_T_66[15:8] ? 8'h6 : _GEN_8356; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8358 = 8'ha6 == _t_T_66[15:8] ? 8'h24 : _GEN_8357; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8359 = 8'ha7 == _t_T_66[15:8] ? 8'h5c : _GEN_8358; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8360 = 8'ha8 == _t_T_66[15:8] ? 8'hc2 : _GEN_8359; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8361 = 8'ha9 == _t_T_66[15:8] ? 8'hd3 : _GEN_8360; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8362 = 8'haa == _t_T_66[15:8] ? 8'hac : _GEN_8361; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8363 = 8'hab == _t_T_66[15:8] ? 8'h62 : _GEN_8362; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8364 = 8'hac == _t_T_66[15:8] ? 8'h91 : _GEN_8363; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8365 = 8'had == _t_T_66[15:8] ? 8'h95 : _GEN_8364; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8366 = 8'hae == _t_T_66[15:8] ? 8'he4 : _GEN_8365; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8367 = 8'haf == _t_T_66[15:8] ? 8'h79 : _GEN_8366; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8368 = 8'hb0 == _t_T_66[15:8] ? 8'he7 : _GEN_8367; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8369 = 8'hb1 == _t_T_66[15:8] ? 8'hc8 : _GEN_8368; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8370 = 8'hb2 == _t_T_66[15:8] ? 8'h37 : _GEN_8369; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8371 = 8'hb3 == _t_T_66[15:8] ? 8'h6d : _GEN_8370; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8372 = 8'hb4 == _t_T_66[15:8] ? 8'h8d : _GEN_8371; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8373 = 8'hb5 == _t_T_66[15:8] ? 8'hd5 : _GEN_8372; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8374 = 8'hb6 == _t_T_66[15:8] ? 8'h4e : _GEN_8373; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8375 = 8'hb7 == _t_T_66[15:8] ? 8'ha9 : _GEN_8374; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8376 = 8'hb8 == _t_T_66[15:8] ? 8'h6c : _GEN_8375; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8377 = 8'hb9 == _t_T_66[15:8] ? 8'h56 : _GEN_8376; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8378 = 8'hba == _t_T_66[15:8] ? 8'hf4 : _GEN_8377; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8379 = 8'hbb == _t_T_66[15:8] ? 8'hea : _GEN_8378; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8380 = 8'hbc == _t_T_66[15:8] ? 8'h65 : _GEN_8379; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8381 = 8'hbd == _t_T_66[15:8] ? 8'h7a : _GEN_8380; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8382 = 8'hbe == _t_T_66[15:8] ? 8'hae : _GEN_8381; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8383 = 8'hbf == _t_T_66[15:8] ? 8'h8 : _GEN_8382; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8384 = 8'hc0 == _t_T_66[15:8] ? 8'hba : _GEN_8383; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8385 = 8'hc1 == _t_T_66[15:8] ? 8'h78 : _GEN_8384; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8386 = 8'hc2 == _t_T_66[15:8] ? 8'h25 : _GEN_8385; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8387 = 8'hc3 == _t_T_66[15:8] ? 8'h2e : _GEN_8386; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8388 = 8'hc4 == _t_T_66[15:8] ? 8'h1c : _GEN_8387; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8389 = 8'hc5 == _t_T_66[15:8] ? 8'ha6 : _GEN_8388; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8390 = 8'hc6 == _t_T_66[15:8] ? 8'hb4 : _GEN_8389; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8391 = 8'hc7 == _t_T_66[15:8] ? 8'hc6 : _GEN_8390; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8392 = 8'hc8 == _t_T_66[15:8] ? 8'he8 : _GEN_8391; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8393 = 8'hc9 == _t_T_66[15:8] ? 8'hdd : _GEN_8392; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8394 = 8'hca == _t_T_66[15:8] ? 8'h74 : _GEN_8393; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8395 = 8'hcb == _t_T_66[15:8] ? 8'h1f : _GEN_8394; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8396 = 8'hcc == _t_T_66[15:8] ? 8'h4b : _GEN_8395; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8397 = 8'hcd == _t_T_66[15:8] ? 8'hbd : _GEN_8396; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8398 = 8'hce == _t_T_66[15:8] ? 8'h8b : _GEN_8397; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8399 = 8'hcf == _t_T_66[15:8] ? 8'h8a : _GEN_8398; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8400 = 8'hd0 == _t_T_66[15:8] ? 8'h70 : _GEN_8399; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8401 = 8'hd1 == _t_T_66[15:8] ? 8'h3e : _GEN_8400; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8402 = 8'hd2 == _t_T_66[15:8] ? 8'hb5 : _GEN_8401; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8403 = 8'hd3 == _t_T_66[15:8] ? 8'h66 : _GEN_8402; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8404 = 8'hd4 == _t_T_66[15:8] ? 8'h48 : _GEN_8403; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8405 = 8'hd5 == _t_T_66[15:8] ? 8'h3 : _GEN_8404; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8406 = 8'hd6 == _t_T_66[15:8] ? 8'hf6 : _GEN_8405; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8407 = 8'hd7 == _t_T_66[15:8] ? 8'he : _GEN_8406; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8408 = 8'hd8 == _t_T_66[15:8] ? 8'h61 : _GEN_8407; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8409 = 8'hd9 == _t_T_66[15:8] ? 8'h35 : _GEN_8408; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8410 = 8'hda == _t_T_66[15:8] ? 8'h57 : _GEN_8409; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8411 = 8'hdb == _t_T_66[15:8] ? 8'hb9 : _GEN_8410; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8412 = 8'hdc == _t_T_66[15:8] ? 8'h86 : _GEN_8411; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8413 = 8'hdd == _t_T_66[15:8] ? 8'hc1 : _GEN_8412; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8414 = 8'hde == _t_T_66[15:8] ? 8'h1d : _GEN_8413; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8415 = 8'hdf == _t_T_66[15:8] ? 8'h9e : _GEN_8414; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8416 = 8'he0 == _t_T_66[15:8] ? 8'he1 : _GEN_8415; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8417 = 8'he1 == _t_T_66[15:8] ? 8'hf8 : _GEN_8416; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8418 = 8'he2 == _t_T_66[15:8] ? 8'h98 : _GEN_8417; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8419 = 8'he3 == _t_T_66[15:8] ? 8'h11 : _GEN_8418; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8420 = 8'he4 == _t_T_66[15:8] ? 8'h69 : _GEN_8419; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8421 = 8'he5 == _t_T_66[15:8] ? 8'hd9 : _GEN_8420; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8422 = 8'he6 == _t_T_66[15:8] ? 8'h8e : _GEN_8421; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8423 = 8'he7 == _t_T_66[15:8] ? 8'h94 : _GEN_8422; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8424 = 8'he8 == _t_T_66[15:8] ? 8'h9b : _GEN_8423; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8425 = 8'he9 == _t_T_66[15:8] ? 8'h1e : _GEN_8424; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8426 = 8'hea == _t_T_66[15:8] ? 8'h87 : _GEN_8425; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8427 = 8'heb == _t_T_66[15:8] ? 8'he9 : _GEN_8426; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8428 = 8'hec == _t_T_66[15:8] ? 8'hce : _GEN_8427; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8429 = 8'hed == _t_T_66[15:8] ? 8'h55 : _GEN_8428; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8430 = 8'hee == _t_T_66[15:8] ? 8'h28 : _GEN_8429; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8431 = 8'hef == _t_T_66[15:8] ? 8'hdf : _GEN_8430; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8432 = 8'hf0 == _t_T_66[15:8] ? 8'h8c : _GEN_8431; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8433 = 8'hf1 == _t_T_66[15:8] ? 8'ha1 : _GEN_8432; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8434 = 8'hf2 == _t_T_66[15:8] ? 8'h89 : _GEN_8433; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8435 = 8'hf3 == _t_T_66[15:8] ? 8'hd : _GEN_8434; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8436 = 8'hf4 == _t_T_66[15:8] ? 8'hbf : _GEN_8435; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8437 = 8'hf5 == _t_T_66[15:8] ? 8'he6 : _GEN_8436; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8438 = 8'hf6 == _t_T_66[15:8] ? 8'h42 : _GEN_8437; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8439 = 8'hf7 == _t_T_66[15:8] ? 8'h68 : _GEN_8438; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8440 = 8'hf8 == _t_T_66[15:8] ? 8'h41 : _GEN_8439; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8441 = 8'hf9 == _t_T_66[15:8] ? 8'h99 : _GEN_8440; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8442 = 8'hfa == _t_T_66[15:8] ? 8'h2d : _GEN_8441; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8443 = 8'hfb == _t_T_66[15:8] ? 8'hf : _GEN_8442; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8444 = 8'hfc == _t_T_66[15:8] ? 8'hb0 : _GEN_8443; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8445 = 8'hfd == _t_T_66[15:8] ? 8'h54 : _GEN_8444; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8446 = 8'hfe == _t_T_66[15:8] ? 8'hbb : _GEN_8445; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8447 = 8'hff == _t_T_66[15:8] ? 8'h16 : _GEN_8446; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8449 = 8'h1 == _t_T_66[7:0] ? 8'h7c : 8'h63; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8450 = 8'h2 == _t_T_66[7:0] ? 8'h77 : _GEN_8449; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8451 = 8'h3 == _t_T_66[7:0] ? 8'h7b : _GEN_8450; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8452 = 8'h4 == _t_T_66[7:0] ? 8'hf2 : _GEN_8451; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8453 = 8'h5 == _t_T_66[7:0] ? 8'h6b : _GEN_8452; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8454 = 8'h6 == _t_T_66[7:0] ? 8'h6f : _GEN_8453; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8455 = 8'h7 == _t_T_66[7:0] ? 8'hc5 : _GEN_8454; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8456 = 8'h8 == _t_T_66[7:0] ? 8'h30 : _GEN_8455; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8457 = 8'h9 == _t_T_66[7:0] ? 8'h1 : _GEN_8456; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8458 = 8'ha == _t_T_66[7:0] ? 8'h67 : _GEN_8457; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8459 = 8'hb == _t_T_66[7:0] ? 8'h2b : _GEN_8458; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8460 = 8'hc == _t_T_66[7:0] ? 8'hfe : _GEN_8459; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8461 = 8'hd == _t_T_66[7:0] ? 8'hd7 : _GEN_8460; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8462 = 8'he == _t_T_66[7:0] ? 8'hab : _GEN_8461; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8463 = 8'hf == _t_T_66[7:0] ? 8'h76 : _GEN_8462; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8464 = 8'h10 == _t_T_66[7:0] ? 8'hca : _GEN_8463; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8465 = 8'h11 == _t_T_66[7:0] ? 8'h82 : _GEN_8464; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8466 = 8'h12 == _t_T_66[7:0] ? 8'hc9 : _GEN_8465; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8467 = 8'h13 == _t_T_66[7:0] ? 8'h7d : _GEN_8466; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8468 = 8'h14 == _t_T_66[7:0] ? 8'hfa : _GEN_8467; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8469 = 8'h15 == _t_T_66[7:0] ? 8'h59 : _GEN_8468; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8470 = 8'h16 == _t_T_66[7:0] ? 8'h47 : _GEN_8469; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8471 = 8'h17 == _t_T_66[7:0] ? 8'hf0 : _GEN_8470; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8472 = 8'h18 == _t_T_66[7:0] ? 8'had : _GEN_8471; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8473 = 8'h19 == _t_T_66[7:0] ? 8'hd4 : _GEN_8472; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8474 = 8'h1a == _t_T_66[7:0] ? 8'ha2 : _GEN_8473; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8475 = 8'h1b == _t_T_66[7:0] ? 8'haf : _GEN_8474; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8476 = 8'h1c == _t_T_66[7:0] ? 8'h9c : _GEN_8475; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8477 = 8'h1d == _t_T_66[7:0] ? 8'ha4 : _GEN_8476; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8478 = 8'h1e == _t_T_66[7:0] ? 8'h72 : _GEN_8477; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8479 = 8'h1f == _t_T_66[7:0] ? 8'hc0 : _GEN_8478; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8480 = 8'h20 == _t_T_66[7:0] ? 8'hb7 : _GEN_8479; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8481 = 8'h21 == _t_T_66[7:0] ? 8'hfd : _GEN_8480; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8482 = 8'h22 == _t_T_66[7:0] ? 8'h93 : _GEN_8481; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8483 = 8'h23 == _t_T_66[7:0] ? 8'h26 : _GEN_8482; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8484 = 8'h24 == _t_T_66[7:0] ? 8'h36 : _GEN_8483; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8485 = 8'h25 == _t_T_66[7:0] ? 8'h3f : _GEN_8484; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8486 = 8'h26 == _t_T_66[7:0] ? 8'hf7 : _GEN_8485; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8487 = 8'h27 == _t_T_66[7:0] ? 8'hcc : _GEN_8486; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8488 = 8'h28 == _t_T_66[7:0] ? 8'h34 : _GEN_8487; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8489 = 8'h29 == _t_T_66[7:0] ? 8'ha5 : _GEN_8488; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8490 = 8'h2a == _t_T_66[7:0] ? 8'he5 : _GEN_8489; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8491 = 8'h2b == _t_T_66[7:0] ? 8'hf1 : _GEN_8490; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8492 = 8'h2c == _t_T_66[7:0] ? 8'h71 : _GEN_8491; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8493 = 8'h2d == _t_T_66[7:0] ? 8'hd8 : _GEN_8492; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8494 = 8'h2e == _t_T_66[7:0] ? 8'h31 : _GEN_8493; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8495 = 8'h2f == _t_T_66[7:0] ? 8'h15 : _GEN_8494; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8496 = 8'h30 == _t_T_66[7:0] ? 8'h4 : _GEN_8495; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8497 = 8'h31 == _t_T_66[7:0] ? 8'hc7 : _GEN_8496; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8498 = 8'h32 == _t_T_66[7:0] ? 8'h23 : _GEN_8497; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8499 = 8'h33 == _t_T_66[7:0] ? 8'hc3 : _GEN_8498; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8500 = 8'h34 == _t_T_66[7:0] ? 8'h18 : _GEN_8499; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8501 = 8'h35 == _t_T_66[7:0] ? 8'h96 : _GEN_8500; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8502 = 8'h36 == _t_T_66[7:0] ? 8'h5 : _GEN_8501; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8503 = 8'h37 == _t_T_66[7:0] ? 8'h9a : _GEN_8502; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8504 = 8'h38 == _t_T_66[7:0] ? 8'h7 : _GEN_8503; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8505 = 8'h39 == _t_T_66[7:0] ? 8'h12 : _GEN_8504; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8506 = 8'h3a == _t_T_66[7:0] ? 8'h80 : _GEN_8505; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8507 = 8'h3b == _t_T_66[7:0] ? 8'he2 : _GEN_8506; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8508 = 8'h3c == _t_T_66[7:0] ? 8'heb : _GEN_8507; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8509 = 8'h3d == _t_T_66[7:0] ? 8'h27 : _GEN_8508; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8510 = 8'h3e == _t_T_66[7:0] ? 8'hb2 : _GEN_8509; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8511 = 8'h3f == _t_T_66[7:0] ? 8'h75 : _GEN_8510; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8512 = 8'h40 == _t_T_66[7:0] ? 8'h9 : _GEN_8511; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8513 = 8'h41 == _t_T_66[7:0] ? 8'h83 : _GEN_8512; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8514 = 8'h42 == _t_T_66[7:0] ? 8'h2c : _GEN_8513; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8515 = 8'h43 == _t_T_66[7:0] ? 8'h1a : _GEN_8514; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8516 = 8'h44 == _t_T_66[7:0] ? 8'h1b : _GEN_8515; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8517 = 8'h45 == _t_T_66[7:0] ? 8'h6e : _GEN_8516; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8518 = 8'h46 == _t_T_66[7:0] ? 8'h5a : _GEN_8517; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8519 = 8'h47 == _t_T_66[7:0] ? 8'ha0 : _GEN_8518; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8520 = 8'h48 == _t_T_66[7:0] ? 8'h52 : _GEN_8519; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8521 = 8'h49 == _t_T_66[7:0] ? 8'h3b : _GEN_8520; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8522 = 8'h4a == _t_T_66[7:0] ? 8'hd6 : _GEN_8521; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8523 = 8'h4b == _t_T_66[7:0] ? 8'hb3 : _GEN_8522; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8524 = 8'h4c == _t_T_66[7:0] ? 8'h29 : _GEN_8523; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8525 = 8'h4d == _t_T_66[7:0] ? 8'he3 : _GEN_8524; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8526 = 8'h4e == _t_T_66[7:0] ? 8'h2f : _GEN_8525; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8527 = 8'h4f == _t_T_66[7:0] ? 8'h84 : _GEN_8526; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8528 = 8'h50 == _t_T_66[7:0] ? 8'h53 : _GEN_8527; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8529 = 8'h51 == _t_T_66[7:0] ? 8'hd1 : _GEN_8528; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8530 = 8'h52 == _t_T_66[7:0] ? 8'h0 : _GEN_8529; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8531 = 8'h53 == _t_T_66[7:0] ? 8'hed : _GEN_8530; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8532 = 8'h54 == _t_T_66[7:0] ? 8'h20 : _GEN_8531; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8533 = 8'h55 == _t_T_66[7:0] ? 8'hfc : _GEN_8532; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8534 = 8'h56 == _t_T_66[7:0] ? 8'hb1 : _GEN_8533; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8535 = 8'h57 == _t_T_66[7:0] ? 8'h5b : _GEN_8534; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8536 = 8'h58 == _t_T_66[7:0] ? 8'h6a : _GEN_8535; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8537 = 8'h59 == _t_T_66[7:0] ? 8'hcb : _GEN_8536; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8538 = 8'h5a == _t_T_66[7:0] ? 8'hbe : _GEN_8537; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8539 = 8'h5b == _t_T_66[7:0] ? 8'h39 : _GEN_8538; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8540 = 8'h5c == _t_T_66[7:0] ? 8'h4a : _GEN_8539; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8541 = 8'h5d == _t_T_66[7:0] ? 8'h4c : _GEN_8540; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8542 = 8'h5e == _t_T_66[7:0] ? 8'h58 : _GEN_8541; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8543 = 8'h5f == _t_T_66[7:0] ? 8'hcf : _GEN_8542; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8544 = 8'h60 == _t_T_66[7:0] ? 8'hd0 : _GEN_8543; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8545 = 8'h61 == _t_T_66[7:0] ? 8'hef : _GEN_8544; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8546 = 8'h62 == _t_T_66[7:0] ? 8'haa : _GEN_8545; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8547 = 8'h63 == _t_T_66[7:0] ? 8'hfb : _GEN_8546; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8548 = 8'h64 == _t_T_66[7:0] ? 8'h43 : _GEN_8547; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8549 = 8'h65 == _t_T_66[7:0] ? 8'h4d : _GEN_8548; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8550 = 8'h66 == _t_T_66[7:0] ? 8'h33 : _GEN_8549; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8551 = 8'h67 == _t_T_66[7:0] ? 8'h85 : _GEN_8550; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8552 = 8'h68 == _t_T_66[7:0] ? 8'h45 : _GEN_8551; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8553 = 8'h69 == _t_T_66[7:0] ? 8'hf9 : _GEN_8552; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8554 = 8'h6a == _t_T_66[7:0] ? 8'h2 : _GEN_8553; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8555 = 8'h6b == _t_T_66[7:0] ? 8'h7f : _GEN_8554; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8556 = 8'h6c == _t_T_66[7:0] ? 8'h50 : _GEN_8555; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8557 = 8'h6d == _t_T_66[7:0] ? 8'h3c : _GEN_8556; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8558 = 8'h6e == _t_T_66[7:0] ? 8'h9f : _GEN_8557; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8559 = 8'h6f == _t_T_66[7:0] ? 8'ha8 : _GEN_8558; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8560 = 8'h70 == _t_T_66[7:0] ? 8'h51 : _GEN_8559; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8561 = 8'h71 == _t_T_66[7:0] ? 8'ha3 : _GEN_8560; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8562 = 8'h72 == _t_T_66[7:0] ? 8'h40 : _GEN_8561; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8563 = 8'h73 == _t_T_66[7:0] ? 8'h8f : _GEN_8562; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8564 = 8'h74 == _t_T_66[7:0] ? 8'h92 : _GEN_8563; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8565 = 8'h75 == _t_T_66[7:0] ? 8'h9d : _GEN_8564; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8566 = 8'h76 == _t_T_66[7:0] ? 8'h38 : _GEN_8565; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8567 = 8'h77 == _t_T_66[7:0] ? 8'hf5 : _GEN_8566; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8568 = 8'h78 == _t_T_66[7:0] ? 8'hbc : _GEN_8567; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8569 = 8'h79 == _t_T_66[7:0] ? 8'hb6 : _GEN_8568; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8570 = 8'h7a == _t_T_66[7:0] ? 8'hda : _GEN_8569; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8571 = 8'h7b == _t_T_66[7:0] ? 8'h21 : _GEN_8570; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8572 = 8'h7c == _t_T_66[7:0] ? 8'h10 : _GEN_8571; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8573 = 8'h7d == _t_T_66[7:0] ? 8'hff : _GEN_8572; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8574 = 8'h7e == _t_T_66[7:0] ? 8'hf3 : _GEN_8573; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8575 = 8'h7f == _t_T_66[7:0] ? 8'hd2 : _GEN_8574; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8576 = 8'h80 == _t_T_66[7:0] ? 8'hcd : _GEN_8575; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8577 = 8'h81 == _t_T_66[7:0] ? 8'hc : _GEN_8576; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8578 = 8'h82 == _t_T_66[7:0] ? 8'h13 : _GEN_8577; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8579 = 8'h83 == _t_T_66[7:0] ? 8'hec : _GEN_8578; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8580 = 8'h84 == _t_T_66[7:0] ? 8'h5f : _GEN_8579; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8581 = 8'h85 == _t_T_66[7:0] ? 8'h97 : _GEN_8580; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8582 = 8'h86 == _t_T_66[7:0] ? 8'h44 : _GEN_8581; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8583 = 8'h87 == _t_T_66[7:0] ? 8'h17 : _GEN_8582; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8584 = 8'h88 == _t_T_66[7:0] ? 8'hc4 : _GEN_8583; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8585 = 8'h89 == _t_T_66[7:0] ? 8'ha7 : _GEN_8584; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8586 = 8'h8a == _t_T_66[7:0] ? 8'h7e : _GEN_8585; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8587 = 8'h8b == _t_T_66[7:0] ? 8'h3d : _GEN_8586; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8588 = 8'h8c == _t_T_66[7:0] ? 8'h64 : _GEN_8587; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8589 = 8'h8d == _t_T_66[7:0] ? 8'h5d : _GEN_8588; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8590 = 8'h8e == _t_T_66[7:0] ? 8'h19 : _GEN_8589; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8591 = 8'h8f == _t_T_66[7:0] ? 8'h73 : _GEN_8590; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8592 = 8'h90 == _t_T_66[7:0] ? 8'h60 : _GEN_8591; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8593 = 8'h91 == _t_T_66[7:0] ? 8'h81 : _GEN_8592; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8594 = 8'h92 == _t_T_66[7:0] ? 8'h4f : _GEN_8593; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8595 = 8'h93 == _t_T_66[7:0] ? 8'hdc : _GEN_8594; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8596 = 8'h94 == _t_T_66[7:0] ? 8'h22 : _GEN_8595; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8597 = 8'h95 == _t_T_66[7:0] ? 8'h2a : _GEN_8596; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8598 = 8'h96 == _t_T_66[7:0] ? 8'h90 : _GEN_8597; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8599 = 8'h97 == _t_T_66[7:0] ? 8'h88 : _GEN_8598; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8600 = 8'h98 == _t_T_66[7:0] ? 8'h46 : _GEN_8599; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8601 = 8'h99 == _t_T_66[7:0] ? 8'hee : _GEN_8600; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8602 = 8'h9a == _t_T_66[7:0] ? 8'hb8 : _GEN_8601; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8603 = 8'h9b == _t_T_66[7:0] ? 8'h14 : _GEN_8602; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8604 = 8'h9c == _t_T_66[7:0] ? 8'hde : _GEN_8603; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8605 = 8'h9d == _t_T_66[7:0] ? 8'h5e : _GEN_8604; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8606 = 8'h9e == _t_T_66[7:0] ? 8'hb : _GEN_8605; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8607 = 8'h9f == _t_T_66[7:0] ? 8'hdb : _GEN_8606; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8608 = 8'ha0 == _t_T_66[7:0] ? 8'he0 : _GEN_8607; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8609 = 8'ha1 == _t_T_66[7:0] ? 8'h32 : _GEN_8608; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8610 = 8'ha2 == _t_T_66[7:0] ? 8'h3a : _GEN_8609; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8611 = 8'ha3 == _t_T_66[7:0] ? 8'ha : _GEN_8610; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8612 = 8'ha4 == _t_T_66[7:0] ? 8'h49 : _GEN_8611; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8613 = 8'ha5 == _t_T_66[7:0] ? 8'h6 : _GEN_8612; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8614 = 8'ha6 == _t_T_66[7:0] ? 8'h24 : _GEN_8613; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8615 = 8'ha7 == _t_T_66[7:0] ? 8'h5c : _GEN_8614; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8616 = 8'ha8 == _t_T_66[7:0] ? 8'hc2 : _GEN_8615; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8617 = 8'ha9 == _t_T_66[7:0] ? 8'hd3 : _GEN_8616; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8618 = 8'haa == _t_T_66[7:0] ? 8'hac : _GEN_8617; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8619 = 8'hab == _t_T_66[7:0] ? 8'h62 : _GEN_8618; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8620 = 8'hac == _t_T_66[7:0] ? 8'h91 : _GEN_8619; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8621 = 8'had == _t_T_66[7:0] ? 8'h95 : _GEN_8620; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8622 = 8'hae == _t_T_66[7:0] ? 8'he4 : _GEN_8621; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8623 = 8'haf == _t_T_66[7:0] ? 8'h79 : _GEN_8622; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8624 = 8'hb0 == _t_T_66[7:0] ? 8'he7 : _GEN_8623; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8625 = 8'hb1 == _t_T_66[7:0] ? 8'hc8 : _GEN_8624; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8626 = 8'hb2 == _t_T_66[7:0] ? 8'h37 : _GEN_8625; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8627 = 8'hb3 == _t_T_66[7:0] ? 8'h6d : _GEN_8626; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8628 = 8'hb4 == _t_T_66[7:0] ? 8'h8d : _GEN_8627; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8629 = 8'hb5 == _t_T_66[7:0] ? 8'hd5 : _GEN_8628; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8630 = 8'hb6 == _t_T_66[7:0] ? 8'h4e : _GEN_8629; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8631 = 8'hb7 == _t_T_66[7:0] ? 8'ha9 : _GEN_8630; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8632 = 8'hb8 == _t_T_66[7:0] ? 8'h6c : _GEN_8631; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8633 = 8'hb9 == _t_T_66[7:0] ? 8'h56 : _GEN_8632; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8634 = 8'hba == _t_T_66[7:0] ? 8'hf4 : _GEN_8633; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8635 = 8'hbb == _t_T_66[7:0] ? 8'hea : _GEN_8634; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8636 = 8'hbc == _t_T_66[7:0] ? 8'h65 : _GEN_8635; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8637 = 8'hbd == _t_T_66[7:0] ? 8'h7a : _GEN_8636; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8638 = 8'hbe == _t_T_66[7:0] ? 8'hae : _GEN_8637; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8639 = 8'hbf == _t_T_66[7:0] ? 8'h8 : _GEN_8638; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8640 = 8'hc0 == _t_T_66[7:0] ? 8'hba : _GEN_8639; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8641 = 8'hc1 == _t_T_66[7:0] ? 8'h78 : _GEN_8640; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8642 = 8'hc2 == _t_T_66[7:0] ? 8'h25 : _GEN_8641; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8643 = 8'hc3 == _t_T_66[7:0] ? 8'h2e : _GEN_8642; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8644 = 8'hc4 == _t_T_66[7:0] ? 8'h1c : _GEN_8643; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8645 = 8'hc5 == _t_T_66[7:0] ? 8'ha6 : _GEN_8644; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8646 = 8'hc6 == _t_T_66[7:0] ? 8'hb4 : _GEN_8645; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8647 = 8'hc7 == _t_T_66[7:0] ? 8'hc6 : _GEN_8646; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8648 = 8'hc8 == _t_T_66[7:0] ? 8'he8 : _GEN_8647; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8649 = 8'hc9 == _t_T_66[7:0] ? 8'hdd : _GEN_8648; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8650 = 8'hca == _t_T_66[7:0] ? 8'h74 : _GEN_8649; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8651 = 8'hcb == _t_T_66[7:0] ? 8'h1f : _GEN_8650; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8652 = 8'hcc == _t_T_66[7:0] ? 8'h4b : _GEN_8651; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8653 = 8'hcd == _t_T_66[7:0] ? 8'hbd : _GEN_8652; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8654 = 8'hce == _t_T_66[7:0] ? 8'h8b : _GEN_8653; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8655 = 8'hcf == _t_T_66[7:0] ? 8'h8a : _GEN_8654; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8656 = 8'hd0 == _t_T_66[7:0] ? 8'h70 : _GEN_8655; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8657 = 8'hd1 == _t_T_66[7:0] ? 8'h3e : _GEN_8656; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8658 = 8'hd2 == _t_T_66[7:0] ? 8'hb5 : _GEN_8657; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8659 = 8'hd3 == _t_T_66[7:0] ? 8'h66 : _GEN_8658; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8660 = 8'hd4 == _t_T_66[7:0] ? 8'h48 : _GEN_8659; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8661 = 8'hd5 == _t_T_66[7:0] ? 8'h3 : _GEN_8660; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8662 = 8'hd6 == _t_T_66[7:0] ? 8'hf6 : _GEN_8661; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8663 = 8'hd7 == _t_T_66[7:0] ? 8'he : _GEN_8662; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8664 = 8'hd8 == _t_T_66[7:0] ? 8'h61 : _GEN_8663; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8665 = 8'hd9 == _t_T_66[7:0] ? 8'h35 : _GEN_8664; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8666 = 8'hda == _t_T_66[7:0] ? 8'h57 : _GEN_8665; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8667 = 8'hdb == _t_T_66[7:0] ? 8'hb9 : _GEN_8666; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8668 = 8'hdc == _t_T_66[7:0] ? 8'h86 : _GEN_8667; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8669 = 8'hdd == _t_T_66[7:0] ? 8'hc1 : _GEN_8668; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8670 = 8'hde == _t_T_66[7:0] ? 8'h1d : _GEN_8669; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8671 = 8'hdf == _t_T_66[7:0] ? 8'h9e : _GEN_8670; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8672 = 8'he0 == _t_T_66[7:0] ? 8'he1 : _GEN_8671; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8673 = 8'he1 == _t_T_66[7:0] ? 8'hf8 : _GEN_8672; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8674 = 8'he2 == _t_T_66[7:0] ? 8'h98 : _GEN_8673; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8675 = 8'he3 == _t_T_66[7:0] ? 8'h11 : _GEN_8674; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8676 = 8'he4 == _t_T_66[7:0] ? 8'h69 : _GEN_8675; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8677 = 8'he5 == _t_T_66[7:0] ? 8'hd9 : _GEN_8676; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8678 = 8'he6 == _t_T_66[7:0] ? 8'h8e : _GEN_8677; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8679 = 8'he7 == _t_T_66[7:0] ? 8'h94 : _GEN_8678; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8680 = 8'he8 == _t_T_66[7:0] ? 8'h9b : _GEN_8679; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8681 = 8'he9 == _t_T_66[7:0] ? 8'h1e : _GEN_8680; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8682 = 8'hea == _t_T_66[7:0] ? 8'h87 : _GEN_8681; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8683 = 8'heb == _t_T_66[7:0] ? 8'he9 : _GEN_8682; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8684 = 8'hec == _t_T_66[7:0] ? 8'hce : _GEN_8683; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8685 = 8'hed == _t_T_66[7:0] ? 8'h55 : _GEN_8684; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8686 = 8'hee == _t_T_66[7:0] ? 8'h28 : _GEN_8685; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8687 = 8'hef == _t_T_66[7:0] ? 8'hdf : _GEN_8686; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8688 = 8'hf0 == _t_T_66[7:0] ? 8'h8c : _GEN_8687; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8689 = 8'hf1 == _t_T_66[7:0] ? 8'ha1 : _GEN_8688; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8690 = 8'hf2 == _t_T_66[7:0] ? 8'h89 : _GEN_8689; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8691 = 8'hf3 == _t_T_66[7:0] ? 8'hd : _GEN_8690; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8692 = 8'hf4 == _t_T_66[7:0] ? 8'hbf : _GEN_8691; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8693 = 8'hf5 == _t_T_66[7:0] ? 8'he6 : _GEN_8692; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8694 = 8'hf6 == _t_T_66[7:0] ? 8'h42 : _GEN_8693; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8695 = 8'hf7 == _t_T_66[7:0] ? 8'h68 : _GEN_8694; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8696 = 8'hf8 == _t_T_66[7:0] ? 8'h41 : _GEN_8695; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8697 = 8'hf9 == _t_T_66[7:0] ? 8'h99 : _GEN_8696; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8698 = 8'hfa == _t_T_66[7:0] ? 8'h2d : _GEN_8697; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8699 = 8'hfb == _t_T_66[7:0] ? 8'hf : _GEN_8698; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8700 = 8'hfc == _t_T_66[7:0] ? 8'hb0 : _GEN_8699; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8701 = 8'hfd == _t_T_66[7:0] ? 8'h54 : _GEN_8700; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8702 = 8'hfe == _t_T_66[7:0] ? 8'hbb : _GEN_8701; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8703 = 8'hff == _t_T_66[7:0] ? 8'h16 : _GEN_8702; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8705 = 8'h1 == _t_T_66[31:24] ? 8'h7c : 8'h63; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8706 = 8'h2 == _t_T_66[31:24] ? 8'h77 : _GEN_8705; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8707 = 8'h3 == _t_T_66[31:24] ? 8'h7b : _GEN_8706; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8708 = 8'h4 == _t_T_66[31:24] ? 8'hf2 : _GEN_8707; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8709 = 8'h5 == _t_T_66[31:24] ? 8'h6b : _GEN_8708; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8710 = 8'h6 == _t_T_66[31:24] ? 8'h6f : _GEN_8709; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8711 = 8'h7 == _t_T_66[31:24] ? 8'hc5 : _GEN_8710; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8712 = 8'h8 == _t_T_66[31:24] ? 8'h30 : _GEN_8711; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8713 = 8'h9 == _t_T_66[31:24] ? 8'h1 : _GEN_8712; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8714 = 8'ha == _t_T_66[31:24] ? 8'h67 : _GEN_8713; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8715 = 8'hb == _t_T_66[31:24] ? 8'h2b : _GEN_8714; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8716 = 8'hc == _t_T_66[31:24] ? 8'hfe : _GEN_8715; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8717 = 8'hd == _t_T_66[31:24] ? 8'hd7 : _GEN_8716; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8718 = 8'he == _t_T_66[31:24] ? 8'hab : _GEN_8717; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8719 = 8'hf == _t_T_66[31:24] ? 8'h76 : _GEN_8718; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8720 = 8'h10 == _t_T_66[31:24] ? 8'hca : _GEN_8719; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8721 = 8'h11 == _t_T_66[31:24] ? 8'h82 : _GEN_8720; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8722 = 8'h12 == _t_T_66[31:24] ? 8'hc9 : _GEN_8721; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8723 = 8'h13 == _t_T_66[31:24] ? 8'h7d : _GEN_8722; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8724 = 8'h14 == _t_T_66[31:24] ? 8'hfa : _GEN_8723; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8725 = 8'h15 == _t_T_66[31:24] ? 8'h59 : _GEN_8724; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8726 = 8'h16 == _t_T_66[31:24] ? 8'h47 : _GEN_8725; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8727 = 8'h17 == _t_T_66[31:24] ? 8'hf0 : _GEN_8726; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8728 = 8'h18 == _t_T_66[31:24] ? 8'had : _GEN_8727; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8729 = 8'h19 == _t_T_66[31:24] ? 8'hd4 : _GEN_8728; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8730 = 8'h1a == _t_T_66[31:24] ? 8'ha2 : _GEN_8729; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8731 = 8'h1b == _t_T_66[31:24] ? 8'haf : _GEN_8730; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8732 = 8'h1c == _t_T_66[31:24] ? 8'h9c : _GEN_8731; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8733 = 8'h1d == _t_T_66[31:24] ? 8'ha4 : _GEN_8732; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8734 = 8'h1e == _t_T_66[31:24] ? 8'h72 : _GEN_8733; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8735 = 8'h1f == _t_T_66[31:24] ? 8'hc0 : _GEN_8734; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8736 = 8'h20 == _t_T_66[31:24] ? 8'hb7 : _GEN_8735; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8737 = 8'h21 == _t_T_66[31:24] ? 8'hfd : _GEN_8736; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8738 = 8'h22 == _t_T_66[31:24] ? 8'h93 : _GEN_8737; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8739 = 8'h23 == _t_T_66[31:24] ? 8'h26 : _GEN_8738; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8740 = 8'h24 == _t_T_66[31:24] ? 8'h36 : _GEN_8739; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8741 = 8'h25 == _t_T_66[31:24] ? 8'h3f : _GEN_8740; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8742 = 8'h26 == _t_T_66[31:24] ? 8'hf7 : _GEN_8741; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8743 = 8'h27 == _t_T_66[31:24] ? 8'hcc : _GEN_8742; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8744 = 8'h28 == _t_T_66[31:24] ? 8'h34 : _GEN_8743; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8745 = 8'h29 == _t_T_66[31:24] ? 8'ha5 : _GEN_8744; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8746 = 8'h2a == _t_T_66[31:24] ? 8'he5 : _GEN_8745; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8747 = 8'h2b == _t_T_66[31:24] ? 8'hf1 : _GEN_8746; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8748 = 8'h2c == _t_T_66[31:24] ? 8'h71 : _GEN_8747; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8749 = 8'h2d == _t_T_66[31:24] ? 8'hd8 : _GEN_8748; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8750 = 8'h2e == _t_T_66[31:24] ? 8'h31 : _GEN_8749; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8751 = 8'h2f == _t_T_66[31:24] ? 8'h15 : _GEN_8750; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8752 = 8'h30 == _t_T_66[31:24] ? 8'h4 : _GEN_8751; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8753 = 8'h31 == _t_T_66[31:24] ? 8'hc7 : _GEN_8752; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8754 = 8'h32 == _t_T_66[31:24] ? 8'h23 : _GEN_8753; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8755 = 8'h33 == _t_T_66[31:24] ? 8'hc3 : _GEN_8754; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8756 = 8'h34 == _t_T_66[31:24] ? 8'h18 : _GEN_8755; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8757 = 8'h35 == _t_T_66[31:24] ? 8'h96 : _GEN_8756; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8758 = 8'h36 == _t_T_66[31:24] ? 8'h5 : _GEN_8757; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8759 = 8'h37 == _t_T_66[31:24] ? 8'h9a : _GEN_8758; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8760 = 8'h38 == _t_T_66[31:24] ? 8'h7 : _GEN_8759; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8761 = 8'h39 == _t_T_66[31:24] ? 8'h12 : _GEN_8760; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8762 = 8'h3a == _t_T_66[31:24] ? 8'h80 : _GEN_8761; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8763 = 8'h3b == _t_T_66[31:24] ? 8'he2 : _GEN_8762; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8764 = 8'h3c == _t_T_66[31:24] ? 8'heb : _GEN_8763; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8765 = 8'h3d == _t_T_66[31:24] ? 8'h27 : _GEN_8764; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8766 = 8'h3e == _t_T_66[31:24] ? 8'hb2 : _GEN_8765; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8767 = 8'h3f == _t_T_66[31:24] ? 8'h75 : _GEN_8766; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8768 = 8'h40 == _t_T_66[31:24] ? 8'h9 : _GEN_8767; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8769 = 8'h41 == _t_T_66[31:24] ? 8'h83 : _GEN_8768; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8770 = 8'h42 == _t_T_66[31:24] ? 8'h2c : _GEN_8769; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8771 = 8'h43 == _t_T_66[31:24] ? 8'h1a : _GEN_8770; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8772 = 8'h44 == _t_T_66[31:24] ? 8'h1b : _GEN_8771; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8773 = 8'h45 == _t_T_66[31:24] ? 8'h6e : _GEN_8772; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8774 = 8'h46 == _t_T_66[31:24] ? 8'h5a : _GEN_8773; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8775 = 8'h47 == _t_T_66[31:24] ? 8'ha0 : _GEN_8774; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8776 = 8'h48 == _t_T_66[31:24] ? 8'h52 : _GEN_8775; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8777 = 8'h49 == _t_T_66[31:24] ? 8'h3b : _GEN_8776; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8778 = 8'h4a == _t_T_66[31:24] ? 8'hd6 : _GEN_8777; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8779 = 8'h4b == _t_T_66[31:24] ? 8'hb3 : _GEN_8778; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8780 = 8'h4c == _t_T_66[31:24] ? 8'h29 : _GEN_8779; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8781 = 8'h4d == _t_T_66[31:24] ? 8'he3 : _GEN_8780; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8782 = 8'h4e == _t_T_66[31:24] ? 8'h2f : _GEN_8781; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8783 = 8'h4f == _t_T_66[31:24] ? 8'h84 : _GEN_8782; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8784 = 8'h50 == _t_T_66[31:24] ? 8'h53 : _GEN_8783; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8785 = 8'h51 == _t_T_66[31:24] ? 8'hd1 : _GEN_8784; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8786 = 8'h52 == _t_T_66[31:24] ? 8'h0 : _GEN_8785; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8787 = 8'h53 == _t_T_66[31:24] ? 8'hed : _GEN_8786; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8788 = 8'h54 == _t_T_66[31:24] ? 8'h20 : _GEN_8787; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8789 = 8'h55 == _t_T_66[31:24] ? 8'hfc : _GEN_8788; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8790 = 8'h56 == _t_T_66[31:24] ? 8'hb1 : _GEN_8789; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8791 = 8'h57 == _t_T_66[31:24] ? 8'h5b : _GEN_8790; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8792 = 8'h58 == _t_T_66[31:24] ? 8'h6a : _GEN_8791; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8793 = 8'h59 == _t_T_66[31:24] ? 8'hcb : _GEN_8792; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8794 = 8'h5a == _t_T_66[31:24] ? 8'hbe : _GEN_8793; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8795 = 8'h5b == _t_T_66[31:24] ? 8'h39 : _GEN_8794; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8796 = 8'h5c == _t_T_66[31:24] ? 8'h4a : _GEN_8795; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8797 = 8'h5d == _t_T_66[31:24] ? 8'h4c : _GEN_8796; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8798 = 8'h5e == _t_T_66[31:24] ? 8'h58 : _GEN_8797; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8799 = 8'h5f == _t_T_66[31:24] ? 8'hcf : _GEN_8798; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8800 = 8'h60 == _t_T_66[31:24] ? 8'hd0 : _GEN_8799; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8801 = 8'h61 == _t_T_66[31:24] ? 8'hef : _GEN_8800; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8802 = 8'h62 == _t_T_66[31:24] ? 8'haa : _GEN_8801; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8803 = 8'h63 == _t_T_66[31:24] ? 8'hfb : _GEN_8802; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8804 = 8'h64 == _t_T_66[31:24] ? 8'h43 : _GEN_8803; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8805 = 8'h65 == _t_T_66[31:24] ? 8'h4d : _GEN_8804; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8806 = 8'h66 == _t_T_66[31:24] ? 8'h33 : _GEN_8805; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8807 = 8'h67 == _t_T_66[31:24] ? 8'h85 : _GEN_8806; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8808 = 8'h68 == _t_T_66[31:24] ? 8'h45 : _GEN_8807; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8809 = 8'h69 == _t_T_66[31:24] ? 8'hf9 : _GEN_8808; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8810 = 8'h6a == _t_T_66[31:24] ? 8'h2 : _GEN_8809; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8811 = 8'h6b == _t_T_66[31:24] ? 8'h7f : _GEN_8810; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8812 = 8'h6c == _t_T_66[31:24] ? 8'h50 : _GEN_8811; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8813 = 8'h6d == _t_T_66[31:24] ? 8'h3c : _GEN_8812; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8814 = 8'h6e == _t_T_66[31:24] ? 8'h9f : _GEN_8813; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8815 = 8'h6f == _t_T_66[31:24] ? 8'ha8 : _GEN_8814; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8816 = 8'h70 == _t_T_66[31:24] ? 8'h51 : _GEN_8815; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8817 = 8'h71 == _t_T_66[31:24] ? 8'ha3 : _GEN_8816; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8818 = 8'h72 == _t_T_66[31:24] ? 8'h40 : _GEN_8817; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8819 = 8'h73 == _t_T_66[31:24] ? 8'h8f : _GEN_8818; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8820 = 8'h74 == _t_T_66[31:24] ? 8'h92 : _GEN_8819; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8821 = 8'h75 == _t_T_66[31:24] ? 8'h9d : _GEN_8820; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8822 = 8'h76 == _t_T_66[31:24] ? 8'h38 : _GEN_8821; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8823 = 8'h77 == _t_T_66[31:24] ? 8'hf5 : _GEN_8822; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8824 = 8'h78 == _t_T_66[31:24] ? 8'hbc : _GEN_8823; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8825 = 8'h79 == _t_T_66[31:24] ? 8'hb6 : _GEN_8824; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8826 = 8'h7a == _t_T_66[31:24] ? 8'hda : _GEN_8825; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8827 = 8'h7b == _t_T_66[31:24] ? 8'h21 : _GEN_8826; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8828 = 8'h7c == _t_T_66[31:24] ? 8'h10 : _GEN_8827; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8829 = 8'h7d == _t_T_66[31:24] ? 8'hff : _GEN_8828; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8830 = 8'h7e == _t_T_66[31:24] ? 8'hf3 : _GEN_8829; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8831 = 8'h7f == _t_T_66[31:24] ? 8'hd2 : _GEN_8830; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8832 = 8'h80 == _t_T_66[31:24] ? 8'hcd : _GEN_8831; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8833 = 8'h81 == _t_T_66[31:24] ? 8'hc : _GEN_8832; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8834 = 8'h82 == _t_T_66[31:24] ? 8'h13 : _GEN_8833; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8835 = 8'h83 == _t_T_66[31:24] ? 8'hec : _GEN_8834; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8836 = 8'h84 == _t_T_66[31:24] ? 8'h5f : _GEN_8835; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8837 = 8'h85 == _t_T_66[31:24] ? 8'h97 : _GEN_8836; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8838 = 8'h86 == _t_T_66[31:24] ? 8'h44 : _GEN_8837; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8839 = 8'h87 == _t_T_66[31:24] ? 8'h17 : _GEN_8838; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8840 = 8'h88 == _t_T_66[31:24] ? 8'hc4 : _GEN_8839; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8841 = 8'h89 == _t_T_66[31:24] ? 8'ha7 : _GEN_8840; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8842 = 8'h8a == _t_T_66[31:24] ? 8'h7e : _GEN_8841; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8843 = 8'h8b == _t_T_66[31:24] ? 8'h3d : _GEN_8842; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8844 = 8'h8c == _t_T_66[31:24] ? 8'h64 : _GEN_8843; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8845 = 8'h8d == _t_T_66[31:24] ? 8'h5d : _GEN_8844; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8846 = 8'h8e == _t_T_66[31:24] ? 8'h19 : _GEN_8845; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8847 = 8'h8f == _t_T_66[31:24] ? 8'h73 : _GEN_8846; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8848 = 8'h90 == _t_T_66[31:24] ? 8'h60 : _GEN_8847; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8849 = 8'h91 == _t_T_66[31:24] ? 8'h81 : _GEN_8848; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8850 = 8'h92 == _t_T_66[31:24] ? 8'h4f : _GEN_8849; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8851 = 8'h93 == _t_T_66[31:24] ? 8'hdc : _GEN_8850; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8852 = 8'h94 == _t_T_66[31:24] ? 8'h22 : _GEN_8851; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8853 = 8'h95 == _t_T_66[31:24] ? 8'h2a : _GEN_8852; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8854 = 8'h96 == _t_T_66[31:24] ? 8'h90 : _GEN_8853; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8855 = 8'h97 == _t_T_66[31:24] ? 8'h88 : _GEN_8854; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8856 = 8'h98 == _t_T_66[31:24] ? 8'h46 : _GEN_8855; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8857 = 8'h99 == _t_T_66[31:24] ? 8'hee : _GEN_8856; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8858 = 8'h9a == _t_T_66[31:24] ? 8'hb8 : _GEN_8857; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8859 = 8'h9b == _t_T_66[31:24] ? 8'h14 : _GEN_8858; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8860 = 8'h9c == _t_T_66[31:24] ? 8'hde : _GEN_8859; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8861 = 8'h9d == _t_T_66[31:24] ? 8'h5e : _GEN_8860; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8862 = 8'h9e == _t_T_66[31:24] ? 8'hb : _GEN_8861; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8863 = 8'h9f == _t_T_66[31:24] ? 8'hdb : _GEN_8862; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8864 = 8'ha0 == _t_T_66[31:24] ? 8'he0 : _GEN_8863; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8865 = 8'ha1 == _t_T_66[31:24] ? 8'h32 : _GEN_8864; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8866 = 8'ha2 == _t_T_66[31:24] ? 8'h3a : _GEN_8865; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8867 = 8'ha3 == _t_T_66[31:24] ? 8'ha : _GEN_8866; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8868 = 8'ha4 == _t_T_66[31:24] ? 8'h49 : _GEN_8867; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8869 = 8'ha5 == _t_T_66[31:24] ? 8'h6 : _GEN_8868; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8870 = 8'ha6 == _t_T_66[31:24] ? 8'h24 : _GEN_8869; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8871 = 8'ha7 == _t_T_66[31:24] ? 8'h5c : _GEN_8870; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8872 = 8'ha8 == _t_T_66[31:24] ? 8'hc2 : _GEN_8871; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8873 = 8'ha9 == _t_T_66[31:24] ? 8'hd3 : _GEN_8872; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8874 = 8'haa == _t_T_66[31:24] ? 8'hac : _GEN_8873; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8875 = 8'hab == _t_T_66[31:24] ? 8'h62 : _GEN_8874; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8876 = 8'hac == _t_T_66[31:24] ? 8'h91 : _GEN_8875; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8877 = 8'had == _t_T_66[31:24] ? 8'h95 : _GEN_8876; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8878 = 8'hae == _t_T_66[31:24] ? 8'he4 : _GEN_8877; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8879 = 8'haf == _t_T_66[31:24] ? 8'h79 : _GEN_8878; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8880 = 8'hb0 == _t_T_66[31:24] ? 8'he7 : _GEN_8879; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8881 = 8'hb1 == _t_T_66[31:24] ? 8'hc8 : _GEN_8880; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8882 = 8'hb2 == _t_T_66[31:24] ? 8'h37 : _GEN_8881; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8883 = 8'hb3 == _t_T_66[31:24] ? 8'h6d : _GEN_8882; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8884 = 8'hb4 == _t_T_66[31:24] ? 8'h8d : _GEN_8883; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8885 = 8'hb5 == _t_T_66[31:24] ? 8'hd5 : _GEN_8884; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8886 = 8'hb6 == _t_T_66[31:24] ? 8'h4e : _GEN_8885; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8887 = 8'hb7 == _t_T_66[31:24] ? 8'ha9 : _GEN_8886; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8888 = 8'hb8 == _t_T_66[31:24] ? 8'h6c : _GEN_8887; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8889 = 8'hb9 == _t_T_66[31:24] ? 8'h56 : _GEN_8888; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8890 = 8'hba == _t_T_66[31:24] ? 8'hf4 : _GEN_8889; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8891 = 8'hbb == _t_T_66[31:24] ? 8'hea : _GEN_8890; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8892 = 8'hbc == _t_T_66[31:24] ? 8'h65 : _GEN_8891; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8893 = 8'hbd == _t_T_66[31:24] ? 8'h7a : _GEN_8892; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8894 = 8'hbe == _t_T_66[31:24] ? 8'hae : _GEN_8893; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8895 = 8'hbf == _t_T_66[31:24] ? 8'h8 : _GEN_8894; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8896 = 8'hc0 == _t_T_66[31:24] ? 8'hba : _GEN_8895; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8897 = 8'hc1 == _t_T_66[31:24] ? 8'h78 : _GEN_8896; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8898 = 8'hc2 == _t_T_66[31:24] ? 8'h25 : _GEN_8897; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8899 = 8'hc3 == _t_T_66[31:24] ? 8'h2e : _GEN_8898; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8900 = 8'hc4 == _t_T_66[31:24] ? 8'h1c : _GEN_8899; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8901 = 8'hc5 == _t_T_66[31:24] ? 8'ha6 : _GEN_8900; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8902 = 8'hc6 == _t_T_66[31:24] ? 8'hb4 : _GEN_8901; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8903 = 8'hc7 == _t_T_66[31:24] ? 8'hc6 : _GEN_8902; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8904 = 8'hc8 == _t_T_66[31:24] ? 8'he8 : _GEN_8903; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8905 = 8'hc9 == _t_T_66[31:24] ? 8'hdd : _GEN_8904; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8906 = 8'hca == _t_T_66[31:24] ? 8'h74 : _GEN_8905; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8907 = 8'hcb == _t_T_66[31:24] ? 8'h1f : _GEN_8906; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8908 = 8'hcc == _t_T_66[31:24] ? 8'h4b : _GEN_8907; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8909 = 8'hcd == _t_T_66[31:24] ? 8'hbd : _GEN_8908; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8910 = 8'hce == _t_T_66[31:24] ? 8'h8b : _GEN_8909; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8911 = 8'hcf == _t_T_66[31:24] ? 8'h8a : _GEN_8910; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8912 = 8'hd0 == _t_T_66[31:24] ? 8'h70 : _GEN_8911; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8913 = 8'hd1 == _t_T_66[31:24] ? 8'h3e : _GEN_8912; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8914 = 8'hd2 == _t_T_66[31:24] ? 8'hb5 : _GEN_8913; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8915 = 8'hd3 == _t_T_66[31:24] ? 8'h66 : _GEN_8914; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8916 = 8'hd4 == _t_T_66[31:24] ? 8'h48 : _GEN_8915; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8917 = 8'hd5 == _t_T_66[31:24] ? 8'h3 : _GEN_8916; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8918 = 8'hd6 == _t_T_66[31:24] ? 8'hf6 : _GEN_8917; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8919 = 8'hd7 == _t_T_66[31:24] ? 8'he : _GEN_8918; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8920 = 8'hd8 == _t_T_66[31:24] ? 8'h61 : _GEN_8919; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8921 = 8'hd9 == _t_T_66[31:24] ? 8'h35 : _GEN_8920; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8922 = 8'hda == _t_T_66[31:24] ? 8'h57 : _GEN_8921; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8923 = 8'hdb == _t_T_66[31:24] ? 8'hb9 : _GEN_8922; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8924 = 8'hdc == _t_T_66[31:24] ? 8'h86 : _GEN_8923; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8925 = 8'hdd == _t_T_66[31:24] ? 8'hc1 : _GEN_8924; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8926 = 8'hde == _t_T_66[31:24] ? 8'h1d : _GEN_8925; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8927 = 8'hdf == _t_T_66[31:24] ? 8'h9e : _GEN_8926; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8928 = 8'he0 == _t_T_66[31:24] ? 8'he1 : _GEN_8927; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8929 = 8'he1 == _t_T_66[31:24] ? 8'hf8 : _GEN_8928; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8930 = 8'he2 == _t_T_66[31:24] ? 8'h98 : _GEN_8929; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8931 = 8'he3 == _t_T_66[31:24] ? 8'h11 : _GEN_8930; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8932 = 8'he4 == _t_T_66[31:24] ? 8'h69 : _GEN_8931; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8933 = 8'he5 == _t_T_66[31:24] ? 8'hd9 : _GEN_8932; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8934 = 8'he6 == _t_T_66[31:24] ? 8'h8e : _GEN_8933; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8935 = 8'he7 == _t_T_66[31:24] ? 8'h94 : _GEN_8934; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8936 = 8'he8 == _t_T_66[31:24] ? 8'h9b : _GEN_8935; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8937 = 8'he9 == _t_T_66[31:24] ? 8'h1e : _GEN_8936; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8938 = 8'hea == _t_T_66[31:24] ? 8'h87 : _GEN_8937; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8939 = 8'heb == _t_T_66[31:24] ? 8'he9 : _GEN_8938; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8940 = 8'hec == _t_T_66[31:24] ? 8'hce : _GEN_8939; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8941 = 8'hed == _t_T_66[31:24] ? 8'h55 : _GEN_8940; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8942 = 8'hee == _t_T_66[31:24] ? 8'h28 : _GEN_8941; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8943 = 8'hef == _t_T_66[31:24] ? 8'hdf : _GEN_8942; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8944 = 8'hf0 == _t_T_66[31:24] ? 8'h8c : _GEN_8943; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8945 = 8'hf1 == _t_T_66[31:24] ? 8'ha1 : _GEN_8944; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8946 = 8'hf2 == _t_T_66[31:24] ? 8'h89 : _GEN_8945; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8947 = 8'hf3 == _t_T_66[31:24] ? 8'hd : _GEN_8946; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8948 = 8'hf4 == _t_T_66[31:24] ? 8'hbf : _GEN_8947; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8949 = 8'hf5 == _t_T_66[31:24] ? 8'he6 : _GEN_8948; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8950 = 8'hf6 == _t_T_66[31:24] ? 8'h42 : _GEN_8949; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8951 = 8'hf7 == _t_T_66[31:24] ? 8'h68 : _GEN_8950; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8952 = 8'hf8 == _t_T_66[31:24] ? 8'h41 : _GEN_8951; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8953 = 8'hf9 == _t_T_66[31:24] ? 8'h99 : _GEN_8952; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8954 = 8'hfa == _t_T_66[31:24] ? 8'h2d : _GEN_8953; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8955 = 8'hfb == _t_T_66[31:24] ? 8'hf : _GEN_8954; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8956 = 8'hfc == _t_T_66[31:24] ? 8'hb0 : _GEN_8955; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8957 = 8'hfd == _t_T_66[31:24] ? 8'h54 : _GEN_8956; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8958 = 8'hfe == _t_T_66[31:24] ? 8'hbb : _GEN_8957; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8959 = 8'hff == _t_T_66[31:24] ? 8'h16 : _GEN_8958; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8961 = 8'h1 == _t_T_66[23:16] ? 8'h7c : 8'h63; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8962 = 8'h2 == _t_T_66[23:16] ? 8'h77 : _GEN_8961; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8963 = 8'h3 == _t_T_66[23:16] ? 8'h7b : _GEN_8962; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8964 = 8'h4 == _t_T_66[23:16] ? 8'hf2 : _GEN_8963; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8965 = 8'h5 == _t_T_66[23:16] ? 8'h6b : _GEN_8964; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8966 = 8'h6 == _t_T_66[23:16] ? 8'h6f : _GEN_8965; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8967 = 8'h7 == _t_T_66[23:16] ? 8'hc5 : _GEN_8966; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8968 = 8'h8 == _t_T_66[23:16] ? 8'h30 : _GEN_8967; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8969 = 8'h9 == _t_T_66[23:16] ? 8'h1 : _GEN_8968; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8970 = 8'ha == _t_T_66[23:16] ? 8'h67 : _GEN_8969; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8971 = 8'hb == _t_T_66[23:16] ? 8'h2b : _GEN_8970; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8972 = 8'hc == _t_T_66[23:16] ? 8'hfe : _GEN_8971; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8973 = 8'hd == _t_T_66[23:16] ? 8'hd7 : _GEN_8972; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8974 = 8'he == _t_T_66[23:16] ? 8'hab : _GEN_8973; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8975 = 8'hf == _t_T_66[23:16] ? 8'h76 : _GEN_8974; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8976 = 8'h10 == _t_T_66[23:16] ? 8'hca : _GEN_8975; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8977 = 8'h11 == _t_T_66[23:16] ? 8'h82 : _GEN_8976; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8978 = 8'h12 == _t_T_66[23:16] ? 8'hc9 : _GEN_8977; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8979 = 8'h13 == _t_T_66[23:16] ? 8'h7d : _GEN_8978; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8980 = 8'h14 == _t_T_66[23:16] ? 8'hfa : _GEN_8979; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8981 = 8'h15 == _t_T_66[23:16] ? 8'h59 : _GEN_8980; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8982 = 8'h16 == _t_T_66[23:16] ? 8'h47 : _GEN_8981; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8983 = 8'h17 == _t_T_66[23:16] ? 8'hf0 : _GEN_8982; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8984 = 8'h18 == _t_T_66[23:16] ? 8'had : _GEN_8983; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8985 = 8'h19 == _t_T_66[23:16] ? 8'hd4 : _GEN_8984; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8986 = 8'h1a == _t_T_66[23:16] ? 8'ha2 : _GEN_8985; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8987 = 8'h1b == _t_T_66[23:16] ? 8'haf : _GEN_8986; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8988 = 8'h1c == _t_T_66[23:16] ? 8'h9c : _GEN_8987; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8989 = 8'h1d == _t_T_66[23:16] ? 8'ha4 : _GEN_8988; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8990 = 8'h1e == _t_T_66[23:16] ? 8'h72 : _GEN_8989; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8991 = 8'h1f == _t_T_66[23:16] ? 8'hc0 : _GEN_8990; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8992 = 8'h20 == _t_T_66[23:16] ? 8'hb7 : _GEN_8991; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8993 = 8'h21 == _t_T_66[23:16] ? 8'hfd : _GEN_8992; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8994 = 8'h22 == _t_T_66[23:16] ? 8'h93 : _GEN_8993; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8995 = 8'h23 == _t_T_66[23:16] ? 8'h26 : _GEN_8994; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8996 = 8'h24 == _t_T_66[23:16] ? 8'h36 : _GEN_8995; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8997 = 8'h25 == _t_T_66[23:16] ? 8'h3f : _GEN_8996; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8998 = 8'h26 == _t_T_66[23:16] ? 8'hf7 : _GEN_8997; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_8999 = 8'h27 == _t_T_66[23:16] ? 8'hcc : _GEN_8998; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9000 = 8'h28 == _t_T_66[23:16] ? 8'h34 : _GEN_8999; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9001 = 8'h29 == _t_T_66[23:16] ? 8'ha5 : _GEN_9000; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9002 = 8'h2a == _t_T_66[23:16] ? 8'he5 : _GEN_9001; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9003 = 8'h2b == _t_T_66[23:16] ? 8'hf1 : _GEN_9002; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9004 = 8'h2c == _t_T_66[23:16] ? 8'h71 : _GEN_9003; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9005 = 8'h2d == _t_T_66[23:16] ? 8'hd8 : _GEN_9004; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9006 = 8'h2e == _t_T_66[23:16] ? 8'h31 : _GEN_9005; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9007 = 8'h2f == _t_T_66[23:16] ? 8'h15 : _GEN_9006; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9008 = 8'h30 == _t_T_66[23:16] ? 8'h4 : _GEN_9007; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9009 = 8'h31 == _t_T_66[23:16] ? 8'hc7 : _GEN_9008; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9010 = 8'h32 == _t_T_66[23:16] ? 8'h23 : _GEN_9009; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9011 = 8'h33 == _t_T_66[23:16] ? 8'hc3 : _GEN_9010; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9012 = 8'h34 == _t_T_66[23:16] ? 8'h18 : _GEN_9011; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9013 = 8'h35 == _t_T_66[23:16] ? 8'h96 : _GEN_9012; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9014 = 8'h36 == _t_T_66[23:16] ? 8'h5 : _GEN_9013; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9015 = 8'h37 == _t_T_66[23:16] ? 8'h9a : _GEN_9014; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9016 = 8'h38 == _t_T_66[23:16] ? 8'h7 : _GEN_9015; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9017 = 8'h39 == _t_T_66[23:16] ? 8'h12 : _GEN_9016; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9018 = 8'h3a == _t_T_66[23:16] ? 8'h80 : _GEN_9017; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9019 = 8'h3b == _t_T_66[23:16] ? 8'he2 : _GEN_9018; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9020 = 8'h3c == _t_T_66[23:16] ? 8'heb : _GEN_9019; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9021 = 8'h3d == _t_T_66[23:16] ? 8'h27 : _GEN_9020; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9022 = 8'h3e == _t_T_66[23:16] ? 8'hb2 : _GEN_9021; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9023 = 8'h3f == _t_T_66[23:16] ? 8'h75 : _GEN_9022; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9024 = 8'h40 == _t_T_66[23:16] ? 8'h9 : _GEN_9023; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9025 = 8'h41 == _t_T_66[23:16] ? 8'h83 : _GEN_9024; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9026 = 8'h42 == _t_T_66[23:16] ? 8'h2c : _GEN_9025; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9027 = 8'h43 == _t_T_66[23:16] ? 8'h1a : _GEN_9026; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9028 = 8'h44 == _t_T_66[23:16] ? 8'h1b : _GEN_9027; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9029 = 8'h45 == _t_T_66[23:16] ? 8'h6e : _GEN_9028; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9030 = 8'h46 == _t_T_66[23:16] ? 8'h5a : _GEN_9029; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9031 = 8'h47 == _t_T_66[23:16] ? 8'ha0 : _GEN_9030; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9032 = 8'h48 == _t_T_66[23:16] ? 8'h52 : _GEN_9031; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9033 = 8'h49 == _t_T_66[23:16] ? 8'h3b : _GEN_9032; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9034 = 8'h4a == _t_T_66[23:16] ? 8'hd6 : _GEN_9033; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9035 = 8'h4b == _t_T_66[23:16] ? 8'hb3 : _GEN_9034; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9036 = 8'h4c == _t_T_66[23:16] ? 8'h29 : _GEN_9035; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9037 = 8'h4d == _t_T_66[23:16] ? 8'he3 : _GEN_9036; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9038 = 8'h4e == _t_T_66[23:16] ? 8'h2f : _GEN_9037; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9039 = 8'h4f == _t_T_66[23:16] ? 8'h84 : _GEN_9038; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9040 = 8'h50 == _t_T_66[23:16] ? 8'h53 : _GEN_9039; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9041 = 8'h51 == _t_T_66[23:16] ? 8'hd1 : _GEN_9040; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9042 = 8'h52 == _t_T_66[23:16] ? 8'h0 : _GEN_9041; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9043 = 8'h53 == _t_T_66[23:16] ? 8'hed : _GEN_9042; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9044 = 8'h54 == _t_T_66[23:16] ? 8'h20 : _GEN_9043; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9045 = 8'h55 == _t_T_66[23:16] ? 8'hfc : _GEN_9044; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9046 = 8'h56 == _t_T_66[23:16] ? 8'hb1 : _GEN_9045; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9047 = 8'h57 == _t_T_66[23:16] ? 8'h5b : _GEN_9046; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9048 = 8'h58 == _t_T_66[23:16] ? 8'h6a : _GEN_9047; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9049 = 8'h59 == _t_T_66[23:16] ? 8'hcb : _GEN_9048; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9050 = 8'h5a == _t_T_66[23:16] ? 8'hbe : _GEN_9049; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9051 = 8'h5b == _t_T_66[23:16] ? 8'h39 : _GEN_9050; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9052 = 8'h5c == _t_T_66[23:16] ? 8'h4a : _GEN_9051; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9053 = 8'h5d == _t_T_66[23:16] ? 8'h4c : _GEN_9052; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9054 = 8'h5e == _t_T_66[23:16] ? 8'h58 : _GEN_9053; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9055 = 8'h5f == _t_T_66[23:16] ? 8'hcf : _GEN_9054; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9056 = 8'h60 == _t_T_66[23:16] ? 8'hd0 : _GEN_9055; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9057 = 8'h61 == _t_T_66[23:16] ? 8'hef : _GEN_9056; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9058 = 8'h62 == _t_T_66[23:16] ? 8'haa : _GEN_9057; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9059 = 8'h63 == _t_T_66[23:16] ? 8'hfb : _GEN_9058; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9060 = 8'h64 == _t_T_66[23:16] ? 8'h43 : _GEN_9059; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9061 = 8'h65 == _t_T_66[23:16] ? 8'h4d : _GEN_9060; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9062 = 8'h66 == _t_T_66[23:16] ? 8'h33 : _GEN_9061; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9063 = 8'h67 == _t_T_66[23:16] ? 8'h85 : _GEN_9062; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9064 = 8'h68 == _t_T_66[23:16] ? 8'h45 : _GEN_9063; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9065 = 8'h69 == _t_T_66[23:16] ? 8'hf9 : _GEN_9064; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9066 = 8'h6a == _t_T_66[23:16] ? 8'h2 : _GEN_9065; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9067 = 8'h6b == _t_T_66[23:16] ? 8'h7f : _GEN_9066; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9068 = 8'h6c == _t_T_66[23:16] ? 8'h50 : _GEN_9067; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9069 = 8'h6d == _t_T_66[23:16] ? 8'h3c : _GEN_9068; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9070 = 8'h6e == _t_T_66[23:16] ? 8'h9f : _GEN_9069; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9071 = 8'h6f == _t_T_66[23:16] ? 8'ha8 : _GEN_9070; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9072 = 8'h70 == _t_T_66[23:16] ? 8'h51 : _GEN_9071; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9073 = 8'h71 == _t_T_66[23:16] ? 8'ha3 : _GEN_9072; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9074 = 8'h72 == _t_T_66[23:16] ? 8'h40 : _GEN_9073; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9075 = 8'h73 == _t_T_66[23:16] ? 8'h8f : _GEN_9074; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9076 = 8'h74 == _t_T_66[23:16] ? 8'h92 : _GEN_9075; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9077 = 8'h75 == _t_T_66[23:16] ? 8'h9d : _GEN_9076; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9078 = 8'h76 == _t_T_66[23:16] ? 8'h38 : _GEN_9077; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9079 = 8'h77 == _t_T_66[23:16] ? 8'hf5 : _GEN_9078; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9080 = 8'h78 == _t_T_66[23:16] ? 8'hbc : _GEN_9079; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9081 = 8'h79 == _t_T_66[23:16] ? 8'hb6 : _GEN_9080; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9082 = 8'h7a == _t_T_66[23:16] ? 8'hda : _GEN_9081; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9083 = 8'h7b == _t_T_66[23:16] ? 8'h21 : _GEN_9082; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9084 = 8'h7c == _t_T_66[23:16] ? 8'h10 : _GEN_9083; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9085 = 8'h7d == _t_T_66[23:16] ? 8'hff : _GEN_9084; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9086 = 8'h7e == _t_T_66[23:16] ? 8'hf3 : _GEN_9085; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9087 = 8'h7f == _t_T_66[23:16] ? 8'hd2 : _GEN_9086; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9088 = 8'h80 == _t_T_66[23:16] ? 8'hcd : _GEN_9087; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9089 = 8'h81 == _t_T_66[23:16] ? 8'hc : _GEN_9088; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9090 = 8'h82 == _t_T_66[23:16] ? 8'h13 : _GEN_9089; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9091 = 8'h83 == _t_T_66[23:16] ? 8'hec : _GEN_9090; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9092 = 8'h84 == _t_T_66[23:16] ? 8'h5f : _GEN_9091; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9093 = 8'h85 == _t_T_66[23:16] ? 8'h97 : _GEN_9092; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9094 = 8'h86 == _t_T_66[23:16] ? 8'h44 : _GEN_9093; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9095 = 8'h87 == _t_T_66[23:16] ? 8'h17 : _GEN_9094; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9096 = 8'h88 == _t_T_66[23:16] ? 8'hc4 : _GEN_9095; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9097 = 8'h89 == _t_T_66[23:16] ? 8'ha7 : _GEN_9096; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9098 = 8'h8a == _t_T_66[23:16] ? 8'h7e : _GEN_9097; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9099 = 8'h8b == _t_T_66[23:16] ? 8'h3d : _GEN_9098; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9100 = 8'h8c == _t_T_66[23:16] ? 8'h64 : _GEN_9099; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9101 = 8'h8d == _t_T_66[23:16] ? 8'h5d : _GEN_9100; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9102 = 8'h8e == _t_T_66[23:16] ? 8'h19 : _GEN_9101; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9103 = 8'h8f == _t_T_66[23:16] ? 8'h73 : _GEN_9102; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9104 = 8'h90 == _t_T_66[23:16] ? 8'h60 : _GEN_9103; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9105 = 8'h91 == _t_T_66[23:16] ? 8'h81 : _GEN_9104; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9106 = 8'h92 == _t_T_66[23:16] ? 8'h4f : _GEN_9105; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9107 = 8'h93 == _t_T_66[23:16] ? 8'hdc : _GEN_9106; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9108 = 8'h94 == _t_T_66[23:16] ? 8'h22 : _GEN_9107; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9109 = 8'h95 == _t_T_66[23:16] ? 8'h2a : _GEN_9108; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9110 = 8'h96 == _t_T_66[23:16] ? 8'h90 : _GEN_9109; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9111 = 8'h97 == _t_T_66[23:16] ? 8'h88 : _GEN_9110; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9112 = 8'h98 == _t_T_66[23:16] ? 8'h46 : _GEN_9111; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9113 = 8'h99 == _t_T_66[23:16] ? 8'hee : _GEN_9112; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9114 = 8'h9a == _t_T_66[23:16] ? 8'hb8 : _GEN_9113; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9115 = 8'h9b == _t_T_66[23:16] ? 8'h14 : _GEN_9114; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9116 = 8'h9c == _t_T_66[23:16] ? 8'hde : _GEN_9115; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9117 = 8'h9d == _t_T_66[23:16] ? 8'h5e : _GEN_9116; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9118 = 8'h9e == _t_T_66[23:16] ? 8'hb : _GEN_9117; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9119 = 8'h9f == _t_T_66[23:16] ? 8'hdb : _GEN_9118; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9120 = 8'ha0 == _t_T_66[23:16] ? 8'he0 : _GEN_9119; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9121 = 8'ha1 == _t_T_66[23:16] ? 8'h32 : _GEN_9120; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9122 = 8'ha2 == _t_T_66[23:16] ? 8'h3a : _GEN_9121; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9123 = 8'ha3 == _t_T_66[23:16] ? 8'ha : _GEN_9122; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9124 = 8'ha4 == _t_T_66[23:16] ? 8'h49 : _GEN_9123; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9125 = 8'ha5 == _t_T_66[23:16] ? 8'h6 : _GEN_9124; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9126 = 8'ha6 == _t_T_66[23:16] ? 8'h24 : _GEN_9125; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9127 = 8'ha7 == _t_T_66[23:16] ? 8'h5c : _GEN_9126; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9128 = 8'ha8 == _t_T_66[23:16] ? 8'hc2 : _GEN_9127; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9129 = 8'ha9 == _t_T_66[23:16] ? 8'hd3 : _GEN_9128; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9130 = 8'haa == _t_T_66[23:16] ? 8'hac : _GEN_9129; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9131 = 8'hab == _t_T_66[23:16] ? 8'h62 : _GEN_9130; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9132 = 8'hac == _t_T_66[23:16] ? 8'h91 : _GEN_9131; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9133 = 8'had == _t_T_66[23:16] ? 8'h95 : _GEN_9132; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9134 = 8'hae == _t_T_66[23:16] ? 8'he4 : _GEN_9133; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9135 = 8'haf == _t_T_66[23:16] ? 8'h79 : _GEN_9134; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9136 = 8'hb0 == _t_T_66[23:16] ? 8'he7 : _GEN_9135; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9137 = 8'hb1 == _t_T_66[23:16] ? 8'hc8 : _GEN_9136; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9138 = 8'hb2 == _t_T_66[23:16] ? 8'h37 : _GEN_9137; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9139 = 8'hb3 == _t_T_66[23:16] ? 8'h6d : _GEN_9138; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9140 = 8'hb4 == _t_T_66[23:16] ? 8'h8d : _GEN_9139; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9141 = 8'hb5 == _t_T_66[23:16] ? 8'hd5 : _GEN_9140; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9142 = 8'hb6 == _t_T_66[23:16] ? 8'h4e : _GEN_9141; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9143 = 8'hb7 == _t_T_66[23:16] ? 8'ha9 : _GEN_9142; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9144 = 8'hb8 == _t_T_66[23:16] ? 8'h6c : _GEN_9143; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9145 = 8'hb9 == _t_T_66[23:16] ? 8'h56 : _GEN_9144; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9146 = 8'hba == _t_T_66[23:16] ? 8'hf4 : _GEN_9145; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9147 = 8'hbb == _t_T_66[23:16] ? 8'hea : _GEN_9146; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9148 = 8'hbc == _t_T_66[23:16] ? 8'h65 : _GEN_9147; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9149 = 8'hbd == _t_T_66[23:16] ? 8'h7a : _GEN_9148; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9150 = 8'hbe == _t_T_66[23:16] ? 8'hae : _GEN_9149; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9151 = 8'hbf == _t_T_66[23:16] ? 8'h8 : _GEN_9150; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9152 = 8'hc0 == _t_T_66[23:16] ? 8'hba : _GEN_9151; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9153 = 8'hc1 == _t_T_66[23:16] ? 8'h78 : _GEN_9152; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9154 = 8'hc2 == _t_T_66[23:16] ? 8'h25 : _GEN_9153; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9155 = 8'hc3 == _t_T_66[23:16] ? 8'h2e : _GEN_9154; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9156 = 8'hc4 == _t_T_66[23:16] ? 8'h1c : _GEN_9155; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9157 = 8'hc5 == _t_T_66[23:16] ? 8'ha6 : _GEN_9156; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9158 = 8'hc6 == _t_T_66[23:16] ? 8'hb4 : _GEN_9157; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9159 = 8'hc7 == _t_T_66[23:16] ? 8'hc6 : _GEN_9158; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9160 = 8'hc8 == _t_T_66[23:16] ? 8'he8 : _GEN_9159; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9161 = 8'hc9 == _t_T_66[23:16] ? 8'hdd : _GEN_9160; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9162 = 8'hca == _t_T_66[23:16] ? 8'h74 : _GEN_9161; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9163 = 8'hcb == _t_T_66[23:16] ? 8'h1f : _GEN_9162; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9164 = 8'hcc == _t_T_66[23:16] ? 8'h4b : _GEN_9163; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9165 = 8'hcd == _t_T_66[23:16] ? 8'hbd : _GEN_9164; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9166 = 8'hce == _t_T_66[23:16] ? 8'h8b : _GEN_9165; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9167 = 8'hcf == _t_T_66[23:16] ? 8'h8a : _GEN_9166; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9168 = 8'hd0 == _t_T_66[23:16] ? 8'h70 : _GEN_9167; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9169 = 8'hd1 == _t_T_66[23:16] ? 8'h3e : _GEN_9168; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9170 = 8'hd2 == _t_T_66[23:16] ? 8'hb5 : _GEN_9169; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9171 = 8'hd3 == _t_T_66[23:16] ? 8'h66 : _GEN_9170; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9172 = 8'hd4 == _t_T_66[23:16] ? 8'h48 : _GEN_9171; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9173 = 8'hd5 == _t_T_66[23:16] ? 8'h3 : _GEN_9172; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9174 = 8'hd6 == _t_T_66[23:16] ? 8'hf6 : _GEN_9173; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9175 = 8'hd7 == _t_T_66[23:16] ? 8'he : _GEN_9174; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9176 = 8'hd8 == _t_T_66[23:16] ? 8'h61 : _GEN_9175; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9177 = 8'hd9 == _t_T_66[23:16] ? 8'h35 : _GEN_9176; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9178 = 8'hda == _t_T_66[23:16] ? 8'h57 : _GEN_9177; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9179 = 8'hdb == _t_T_66[23:16] ? 8'hb9 : _GEN_9178; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9180 = 8'hdc == _t_T_66[23:16] ? 8'h86 : _GEN_9179; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9181 = 8'hdd == _t_T_66[23:16] ? 8'hc1 : _GEN_9180; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9182 = 8'hde == _t_T_66[23:16] ? 8'h1d : _GEN_9181; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9183 = 8'hdf == _t_T_66[23:16] ? 8'h9e : _GEN_9182; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9184 = 8'he0 == _t_T_66[23:16] ? 8'he1 : _GEN_9183; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9185 = 8'he1 == _t_T_66[23:16] ? 8'hf8 : _GEN_9184; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9186 = 8'he2 == _t_T_66[23:16] ? 8'h98 : _GEN_9185; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9187 = 8'he3 == _t_T_66[23:16] ? 8'h11 : _GEN_9186; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9188 = 8'he4 == _t_T_66[23:16] ? 8'h69 : _GEN_9187; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9189 = 8'he5 == _t_T_66[23:16] ? 8'hd9 : _GEN_9188; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9190 = 8'he6 == _t_T_66[23:16] ? 8'h8e : _GEN_9189; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9191 = 8'he7 == _t_T_66[23:16] ? 8'h94 : _GEN_9190; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9192 = 8'he8 == _t_T_66[23:16] ? 8'h9b : _GEN_9191; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9193 = 8'he9 == _t_T_66[23:16] ? 8'h1e : _GEN_9192; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9194 = 8'hea == _t_T_66[23:16] ? 8'h87 : _GEN_9193; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9195 = 8'heb == _t_T_66[23:16] ? 8'he9 : _GEN_9194; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9196 = 8'hec == _t_T_66[23:16] ? 8'hce : _GEN_9195; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9197 = 8'hed == _t_T_66[23:16] ? 8'h55 : _GEN_9196; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9198 = 8'hee == _t_T_66[23:16] ? 8'h28 : _GEN_9197; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9199 = 8'hef == _t_T_66[23:16] ? 8'hdf : _GEN_9198; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9200 = 8'hf0 == _t_T_66[23:16] ? 8'h8c : _GEN_9199; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9201 = 8'hf1 == _t_T_66[23:16] ? 8'ha1 : _GEN_9200; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9202 = 8'hf2 == _t_T_66[23:16] ? 8'h89 : _GEN_9201; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9203 = 8'hf3 == _t_T_66[23:16] ? 8'hd : _GEN_9202; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9204 = 8'hf4 == _t_T_66[23:16] ? 8'hbf : _GEN_9203; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9205 = 8'hf5 == _t_T_66[23:16] ? 8'he6 : _GEN_9204; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9206 = 8'hf6 == _t_T_66[23:16] ? 8'h42 : _GEN_9205; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9207 = 8'hf7 == _t_T_66[23:16] ? 8'h68 : _GEN_9206; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9208 = 8'hf8 == _t_T_66[23:16] ? 8'h41 : _GEN_9207; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9209 = 8'hf9 == _t_T_66[23:16] ? 8'h99 : _GEN_9208; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9210 = 8'hfa == _t_T_66[23:16] ? 8'h2d : _GEN_9209; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9211 = 8'hfb == _t_T_66[23:16] ? 8'hf : _GEN_9210; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9212 = 8'hfc == _t_T_66[23:16] ? 8'hb0 : _GEN_9211; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9213 = 8'hfd == _t_T_66[23:16] ? 8'h54 : _GEN_9212; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9214 = 8'hfe == _t_T_66[23:16] ? 8'hbb : _GEN_9213; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9215 = 8'hff == _t_T_66[23:16] ? 8'h16 : _GEN_9214; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [31:0] _t_T_71 = {_GEN_8959,_GEN_9215,_GEN_8447,_GEN_8703}; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:8]
  wire [31:0] t_8 = _t_T_71 ^ 32'h1b000000; // @[src/main/scala/crypto/aes/KeySchedule.scala 59:32]
  wire [31:0] w_36 = w_32 ^ t_8; // @[src/main/scala/crypto/aes/KeySchedule.scala 63:21]
  wire [31:0] w_37 = w_33 ^ w_36; // @[src/main/scala/crypto/aes/KeySchedule.scala 63:21]
  wire [31:0] w_38 = w_34 ^ w_37; // @[src/main/scala/crypto/aes/KeySchedule.scala 63:21]
  wire [31:0] w_39 = w_35 ^ w_38; // @[src/main/scala/crypto/aes/KeySchedule.scala 63:21]
  wire [31:0] _t_T_74 = {w_39[23:0],w_39[31:24]}; // @[src/main/scala/crypto/aes/KeySchedule.scala 23:43]
  wire [7:0] _GEN_9217 = 8'h1 == _t_T_74[15:8] ? 8'h7c : 8'h63; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9218 = 8'h2 == _t_T_74[15:8] ? 8'h77 : _GEN_9217; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9219 = 8'h3 == _t_T_74[15:8] ? 8'h7b : _GEN_9218; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9220 = 8'h4 == _t_T_74[15:8] ? 8'hf2 : _GEN_9219; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9221 = 8'h5 == _t_T_74[15:8] ? 8'h6b : _GEN_9220; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9222 = 8'h6 == _t_T_74[15:8] ? 8'h6f : _GEN_9221; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9223 = 8'h7 == _t_T_74[15:8] ? 8'hc5 : _GEN_9222; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9224 = 8'h8 == _t_T_74[15:8] ? 8'h30 : _GEN_9223; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9225 = 8'h9 == _t_T_74[15:8] ? 8'h1 : _GEN_9224; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9226 = 8'ha == _t_T_74[15:8] ? 8'h67 : _GEN_9225; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9227 = 8'hb == _t_T_74[15:8] ? 8'h2b : _GEN_9226; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9228 = 8'hc == _t_T_74[15:8] ? 8'hfe : _GEN_9227; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9229 = 8'hd == _t_T_74[15:8] ? 8'hd7 : _GEN_9228; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9230 = 8'he == _t_T_74[15:8] ? 8'hab : _GEN_9229; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9231 = 8'hf == _t_T_74[15:8] ? 8'h76 : _GEN_9230; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9232 = 8'h10 == _t_T_74[15:8] ? 8'hca : _GEN_9231; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9233 = 8'h11 == _t_T_74[15:8] ? 8'h82 : _GEN_9232; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9234 = 8'h12 == _t_T_74[15:8] ? 8'hc9 : _GEN_9233; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9235 = 8'h13 == _t_T_74[15:8] ? 8'h7d : _GEN_9234; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9236 = 8'h14 == _t_T_74[15:8] ? 8'hfa : _GEN_9235; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9237 = 8'h15 == _t_T_74[15:8] ? 8'h59 : _GEN_9236; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9238 = 8'h16 == _t_T_74[15:8] ? 8'h47 : _GEN_9237; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9239 = 8'h17 == _t_T_74[15:8] ? 8'hf0 : _GEN_9238; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9240 = 8'h18 == _t_T_74[15:8] ? 8'had : _GEN_9239; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9241 = 8'h19 == _t_T_74[15:8] ? 8'hd4 : _GEN_9240; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9242 = 8'h1a == _t_T_74[15:8] ? 8'ha2 : _GEN_9241; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9243 = 8'h1b == _t_T_74[15:8] ? 8'haf : _GEN_9242; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9244 = 8'h1c == _t_T_74[15:8] ? 8'h9c : _GEN_9243; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9245 = 8'h1d == _t_T_74[15:8] ? 8'ha4 : _GEN_9244; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9246 = 8'h1e == _t_T_74[15:8] ? 8'h72 : _GEN_9245; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9247 = 8'h1f == _t_T_74[15:8] ? 8'hc0 : _GEN_9246; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9248 = 8'h20 == _t_T_74[15:8] ? 8'hb7 : _GEN_9247; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9249 = 8'h21 == _t_T_74[15:8] ? 8'hfd : _GEN_9248; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9250 = 8'h22 == _t_T_74[15:8] ? 8'h93 : _GEN_9249; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9251 = 8'h23 == _t_T_74[15:8] ? 8'h26 : _GEN_9250; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9252 = 8'h24 == _t_T_74[15:8] ? 8'h36 : _GEN_9251; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9253 = 8'h25 == _t_T_74[15:8] ? 8'h3f : _GEN_9252; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9254 = 8'h26 == _t_T_74[15:8] ? 8'hf7 : _GEN_9253; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9255 = 8'h27 == _t_T_74[15:8] ? 8'hcc : _GEN_9254; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9256 = 8'h28 == _t_T_74[15:8] ? 8'h34 : _GEN_9255; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9257 = 8'h29 == _t_T_74[15:8] ? 8'ha5 : _GEN_9256; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9258 = 8'h2a == _t_T_74[15:8] ? 8'he5 : _GEN_9257; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9259 = 8'h2b == _t_T_74[15:8] ? 8'hf1 : _GEN_9258; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9260 = 8'h2c == _t_T_74[15:8] ? 8'h71 : _GEN_9259; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9261 = 8'h2d == _t_T_74[15:8] ? 8'hd8 : _GEN_9260; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9262 = 8'h2e == _t_T_74[15:8] ? 8'h31 : _GEN_9261; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9263 = 8'h2f == _t_T_74[15:8] ? 8'h15 : _GEN_9262; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9264 = 8'h30 == _t_T_74[15:8] ? 8'h4 : _GEN_9263; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9265 = 8'h31 == _t_T_74[15:8] ? 8'hc7 : _GEN_9264; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9266 = 8'h32 == _t_T_74[15:8] ? 8'h23 : _GEN_9265; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9267 = 8'h33 == _t_T_74[15:8] ? 8'hc3 : _GEN_9266; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9268 = 8'h34 == _t_T_74[15:8] ? 8'h18 : _GEN_9267; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9269 = 8'h35 == _t_T_74[15:8] ? 8'h96 : _GEN_9268; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9270 = 8'h36 == _t_T_74[15:8] ? 8'h5 : _GEN_9269; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9271 = 8'h37 == _t_T_74[15:8] ? 8'h9a : _GEN_9270; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9272 = 8'h38 == _t_T_74[15:8] ? 8'h7 : _GEN_9271; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9273 = 8'h39 == _t_T_74[15:8] ? 8'h12 : _GEN_9272; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9274 = 8'h3a == _t_T_74[15:8] ? 8'h80 : _GEN_9273; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9275 = 8'h3b == _t_T_74[15:8] ? 8'he2 : _GEN_9274; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9276 = 8'h3c == _t_T_74[15:8] ? 8'heb : _GEN_9275; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9277 = 8'h3d == _t_T_74[15:8] ? 8'h27 : _GEN_9276; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9278 = 8'h3e == _t_T_74[15:8] ? 8'hb2 : _GEN_9277; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9279 = 8'h3f == _t_T_74[15:8] ? 8'h75 : _GEN_9278; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9280 = 8'h40 == _t_T_74[15:8] ? 8'h9 : _GEN_9279; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9281 = 8'h41 == _t_T_74[15:8] ? 8'h83 : _GEN_9280; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9282 = 8'h42 == _t_T_74[15:8] ? 8'h2c : _GEN_9281; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9283 = 8'h43 == _t_T_74[15:8] ? 8'h1a : _GEN_9282; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9284 = 8'h44 == _t_T_74[15:8] ? 8'h1b : _GEN_9283; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9285 = 8'h45 == _t_T_74[15:8] ? 8'h6e : _GEN_9284; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9286 = 8'h46 == _t_T_74[15:8] ? 8'h5a : _GEN_9285; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9287 = 8'h47 == _t_T_74[15:8] ? 8'ha0 : _GEN_9286; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9288 = 8'h48 == _t_T_74[15:8] ? 8'h52 : _GEN_9287; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9289 = 8'h49 == _t_T_74[15:8] ? 8'h3b : _GEN_9288; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9290 = 8'h4a == _t_T_74[15:8] ? 8'hd6 : _GEN_9289; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9291 = 8'h4b == _t_T_74[15:8] ? 8'hb3 : _GEN_9290; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9292 = 8'h4c == _t_T_74[15:8] ? 8'h29 : _GEN_9291; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9293 = 8'h4d == _t_T_74[15:8] ? 8'he3 : _GEN_9292; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9294 = 8'h4e == _t_T_74[15:8] ? 8'h2f : _GEN_9293; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9295 = 8'h4f == _t_T_74[15:8] ? 8'h84 : _GEN_9294; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9296 = 8'h50 == _t_T_74[15:8] ? 8'h53 : _GEN_9295; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9297 = 8'h51 == _t_T_74[15:8] ? 8'hd1 : _GEN_9296; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9298 = 8'h52 == _t_T_74[15:8] ? 8'h0 : _GEN_9297; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9299 = 8'h53 == _t_T_74[15:8] ? 8'hed : _GEN_9298; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9300 = 8'h54 == _t_T_74[15:8] ? 8'h20 : _GEN_9299; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9301 = 8'h55 == _t_T_74[15:8] ? 8'hfc : _GEN_9300; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9302 = 8'h56 == _t_T_74[15:8] ? 8'hb1 : _GEN_9301; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9303 = 8'h57 == _t_T_74[15:8] ? 8'h5b : _GEN_9302; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9304 = 8'h58 == _t_T_74[15:8] ? 8'h6a : _GEN_9303; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9305 = 8'h59 == _t_T_74[15:8] ? 8'hcb : _GEN_9304; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9306 = 8'h5a == _t_T_74[15:8] ? 8'hbe : _GEN_9305; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9307 = 8'h5b == _t_T_74[15:8] ? 8'h39 : _GEN_9306; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9308 = 8'h5c == _t_T_74[15:8] ? 8'h4a : _GEN_9307; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9309 = 8'h5d == _t_T_74[15:8] ? 8'h4c : _GEN_9308; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9310 = 8'h5e == _t_T_74[15:8] ? 8'h58 : _GEN_9309; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9311 = 8'h5f == _t_T_74[15:8] ? 8'hcf : _GEN_9310; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9312 = 8'h60 == _t_T_74[15:8] ? 8'hd0 : _GEN_9311; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9313 = 8'h61 == _t_T_74[15:8] ? 8'hef : _GEN_9312; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9314 = 8'h62 == _t_T_74[15:8] ? 8'haa : _GEN_9313; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9315 = 8'h63 == _t_T_74[15:8] ? 8'hfb : _GEN_9314; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9316 = 8'h64 == _t_T_74[15:8] ? 8'h43 : _GEN_9315; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9317 = 8'h65 == _t_T_74[15:8] ? 8'h4d : _GEN_9316; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9318 = 8'h66 == _t_T_74[15:8] ? 8'h33 : _GEN_9317; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9319 = 8'h67 == _t_T_74[15:8] ? 8'h85 : _GEN_9318; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9320 = 8'h68 == _t_T_74[15:8] ? 8'h45 : _GEN_9319; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9321 = 8'h69 == _t_T_74[15:8] ? 8'hf9 : _GEN_9320; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9322 = 8'h6a == _t_T_74[15:8] ? 8'h2 : _GEN_9321; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9323 = 8'h6b == _t_T_74[15:8] ? 8'h7f : _GEN_9322; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9324 = 8'h6c == _t_T_74[15:8] ? 8'h50 : _GEN_9323; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9325 = 8'h6d == _t_T_74[15:8] ? 8'h3c : _GEN_9324; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9326 = 8'h6e == _t_T_74[15:8] ? 8'h9f : _GEN_9325; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9327 = 8'h6f == _t_T_74[15:8] ? 8'ha8 : _GEN_9326; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9328 = 8'h70 == _t_T_74[15:8] ? 8'h51 : _GEN_9327; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9329 = 8'h71 == _t_T_74[15:8] ? 8'ha3 : _GEN_9328; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9330 = 8'h72 == _t_T_74[15:8] ? 8'h40 : _GEN_9329; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9331 = 8'h73 == _t_T_74[15:8] ? 8'h8f : _GEN_9330; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9332 = 8'h74 == _t_T_74[15:8] ? 8'h92 : _GEN_9331; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9333 = 8'h75 == _t_T_74[15:8] ? 8'h9d : _GEN_9332; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9334 = 8'h76 == _t_T_74[15:8] ? 8'h38 : _GEN_9333; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9335 = 8'h77 == _t_T_74[15:8] ? 8'hf5 : _GEN_9334; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9336 = 8'h78 == _t_T_74[15:8] ? 8'hbc : _GEN_9335; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9337 = 8'h79 == _t_T_74[15:8] ? 8'hb6 : _GEN_9336; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9338 = 8'h7a == _t_T_74[15:8] ? 8'hda : _GEN_9337; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9339 = 8'h7b == _t_T_74[15:8] ? 8'h21 : _GEN_9338; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9340 = 8'h7c == _t_T_74[15:8] ? 8'h10 : _GEN_9339; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9341 = 8'h7d == _t_T_74[15:8] ? 8'hff : _GEN_9340; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9342 = 8'h7e == _t_T_74[15:8] ? 8'hf3 : _GEN_9341; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9343 = 8'h7f == _t_T_74[15:8] ? 8'hd2 : _GEN_9342; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9344 = 8'h80 == _t_T_74[15:8] ? 8'hcd : _GEN_9343; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9345 = 8'h81 == _t_T_74[15:8] ? 8'hc : _GEN_9344; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9346 = 8'h82 == _t_T_74[15:8] ? 8'h13 : _GEN_9345; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9347 = 8'h83 == _t_T_74[15:8] ? 8'hec : _GEN_9346; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9348 = 8'h84 == _t_T_74[15:8] ? 8'h5f : _GEN_9347; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9349 = 8'h85 == _t_T_74[15:8] ? 8'h97 : _GEN_9348; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9350 = 8'h86 == _t_T_74[15:8] ? 8'h44 : _GEN_9349; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9351 = 8'h87 == _t_T_74[15:8] ? 8'h17 : _GEN_9350; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9352 = 8'h88 == _t_T_74[15:8] ? 8'hc4 : _GEN_9351; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9353 = 8'h89 == _t_T_74[15:8] ? 8'ha7 : _GEN_9352; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9354 = 8'h8a == _t_T_74[15:8] ? 8'h7e : _GEN_9353; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9355 = 8'h8b == _t_T_74[15:8] ? 8'h3d : _GEN_9354; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9356 = 8'h8c == _t_T_74[15:8] ? 8'h64 : _GEN_9355; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9357 = 8'h8d == _t_T_74[15:8] ? 8'h5d : _GEN_9356; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9358 = 8'h8e == _t_T_74[15:8] ? 8'h19 : _GEN_9357; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9359 = 8'h8f == _t_T_74[15:8] ? 8'h73 : _GEN_9358; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9360 = 8'h90 == _t_T_74[15:8] ? 8'h60 : _GEN_9359; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9361 = 8'h91 == _t_T_74[15:8] ? 8'h81 : _GEN_9360; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9362 = 8'h92 == _t_T_74[15:8] ? 8'h4f : _GEN_9361; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9363 = 8'h93 == _t_T_74[15:8] ? 8'hdc : _GEN_9362; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9364 = 8'h94 == _t_T_74[15:8] ? 8'h22 : _GEN_9363; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9365 = 8'h95 == _t_T_74[15:8] ? 8'h2a : _GEN_9364; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9366 = 8'h96 == _t_T_74[15:8] ? 8'h90 : _GEN_9365; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9367 = 8'h97 == _t_T_74[15:8] ? 8'h88 : _GEN_9366; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9368 = 8'h98 == _t_T_74[15:8] ? 8'h46 : _GEN_9367; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9369 = 8'h99 == _t_T_74[15:8] ? 8'hee : _GEN_9368; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9370 = 8'h9a == _t_T_74[15:8] ? 8'hb8 : _GEN_9369; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9371 = 8'h9b == _t_T_74[15:8] ? 8'h14 : _GEN_9370; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9372 = 8'h9c == _t_T_74[15:8] ? 8'hde : _GEN_9371; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9373 = 8'h9d == _t_T_74[15:8] ? 8'h5e : _GEN_9372; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9374 = 8'h9e == _t_T_74[15:8] ? 8'hb : _GEN_9373; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9375 = 8'h9f == _t_T_74[15:8] ? 8'hdb : _GEN_9374; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9376 = 8'ha0 == _t_T_74[15:8] ? 8'he0 : _GEN_9375; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9377 = 8'ha1 == _t_T_74[15:8] ? 8'h32 : _GEN_9376; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9378 = 8'ha2 == _t_T_74[15:8] ? 8'h3a : _GEN_9377; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9379 = 8'ha3 == _t_T_74[15:8] ? 8'ha : _GEN_9378; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9380 = 8'ha4 == _t_T_74[15:8] ? 8'h49 : _GEN_9379; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9381 = 8'ha5 == _t_T_74[15:8] ? 8'h6 : _GEN_9380; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9382 = 8'ha6 == _t_T_74[15:8] ? 8'h24 : _GEN_9381; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9383 = 8'ha7 == _t_T_74[15:8] ? 8'h5c : _GEN_9382; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9384 = 8'ha8 == _t_T_74[15:8] ? 8'hc2 : _GEN_9383; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9385 = 8'ha9 == _t_T_74[15:8] ? 8'hd3 : _GEN_9384; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9386 = 8'haa == _t_T_74[15:8] ? 8'hac : _GEN_9385; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9387 = 8'hab == _t_T_74[15:8] ? 8'h62 : _GEN_9386; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9388 = 8'hac == _t_T_74[15:8] ? 8'h91 : _GEN_9387; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9389 = 8'had == _t_T_74[15:8] ? 8'h95 : _GEN_9388; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9390 = 8'hae == _t_T_74[15:8] ? 8'he4 : _GEN_9389; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9391 = 8'haf == _t_T_74[15:8] ? 8'h79 : _GEN_9390; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9392 = 8'hb0 == _t_T_74[15:8] ? 8'he7 : _GEN_9391; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9393 = 8'hb1 == _t_T_74[15:8] ? 8'hc8 : _GEN_9392; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9394 = 8'hb2 == _t_T_74[15:8] ? 8'h37 : _GEN_9393; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9395 = 8'hb3 == _t_T_74[15:8] ? 8'h6d : _GEN_9394; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9396 = 8'hb4 == _t_T_74[15:8] ? 8'h8d : _GEN_9395; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9397 = 8'hb5 == _t_T_74[15:8] ? 8'hd5 : _GEN_9396; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9398 = 8'hb6 == _t_T_74[15:8] ? 8'h4e : _GEN_9397; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9399 = 8'hb7 == _t_T_74[15:8] ? 8'ha9 : _GEN_9398; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9400 = 8'hb8 == _t_T_74[15:8] ? 8'h6c : _GEN_9399; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9401 = 8'hb9 == _t_T_74[15:8] ? 8'h56 : _GEN_9400; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9402 = 8'hba == _t_T_74[15:8] ? 8'hf4 : _GEN_9401; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9403 = 8'hbb == _t_T_74[15:8] ? 8'hea : _GEN_9402; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9404 = 8'hbc == _t_T_74[15:8] ? 8'h65 : _GEN_9403; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9405 = 8'hbd == _t_T_74[15:8] ? 8'h7a : _GEN_9404; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9406 = 8'hbe == _t_T_74[15:8] ? 8'hae : _GEN_9405; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9407 = 8'hbf == _t_T_74[15:8] ? 8'h8 : _GEN_9406; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9408 = 8'hc0 == _t_T_74[15:8] ? 8'hba : _GEN_9407; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9409 = 8'hc1 == _t_T_74[15:8] ? 8'h78 : _GEN_9408; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9410 = 8'hc2 == _t_T_74[15:8] ? 8'h25 : _GEN_9409; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9411 = 8'hc3 == _t_T_74[15:8] ? 8'h2e : _GEN_9410; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9412 = 8'hc4 == _t_T_74[15:8] ? 8'h1c : _GEN_9411; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9413 = 8'hc5 == _t_T_74[15:8] ? 8'ha6 : _GEN_9412; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9414 = 8'hc6 == _t_T_74[15:8] ? 8'hb4 : _GEN_9413; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9415 = 8'hc7 == _t_T_74[15:8] ? 8'hc6 : _GEN_9414; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9416 = 8'hc8 == _t_T_74[15:8] ? 8'he8 : _GEN_9415; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9417 = 8'hc9 == _t_T_74[15:8] ? 8'hdd : _GEN_9416; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9418 = 8'hca == _t_T_74[15:8] ? 8'h74 : _GEN_9417; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9419 = 8'hcb == _t_T_74[15:8] ? 8'h1f : _GEN_9418; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9420 = 8'hcc == _t_T_74[15:8] ? 8'h4b : _GEN_9419; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9421 = 8'hcd == _t_T_74[15:8] ? 8'hbd : _GEN_9420; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9422 = 8'hce == _t_T_74[15:8] ? 8'h8b : _GEN_9421; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9423 = 8'hcf == _t_T_74[15:8] ? 8'h8a : _GEN_9422; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9424 = 8'hd0 == _t_T_74[15:8] ? 8'h70 : _GEN_9423; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9425 = 8'hd1 == _t_T_74[15:8] ? 8'h3e : _GEN_9424; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9426 = 8'hd2 == _t_T_74[15:8] ? 8'hb5 : _GEN_9425; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9427 = 8'hd3 == _t_T_74[15:8] ? 8'h66 : _GEN_9426; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9428 = 8'hd4 == _t_T_74[15:8] ? 8'h48 : _GEN_9427; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9429 = 8'hd5 == _t_T_74[15:8] ? 8'h3 : _GEN_9428; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9430 = 8'hd6 == _t_T_74[15:8] ? 8'hf6 : _GEN_9429; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9431 = 8'hd7 == _t_T_74[15:8] ? 8'he : _GEN_9430; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9432 = 8'hd8 == _t_T_74[15:8] ? 8'h61 : _GEN_9431; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9433 = 8'hd9 == _t_T_74[15:8] ? 8'h35 : _GEN_9432; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9434 = 8'hda == _t_T_74[15:8] ? 8'h57 : _GEN_9433; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9435 = 8'hdb == _t_T_74[15:8] ? 8'hb9 : _GEN_9434; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9436 = 8'hdc == _t_T_74[15:8] ? 8'h86 : _GEN_9435; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9437 = 8'hdd == _t_T_74[15:8] ? 8'hc1 : _GEN_9436; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9438 = 8'hde == _t_T_74[15:8] ? 8'h1d : _GEN_9437; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9439 = 8'hdf == _t_T_74[15:8] ? 8'h9e : _GEN_9438; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9440 = 8'he0 == _t_T_74[15:8] ? 8'he1 : _GEN_9439; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9441 = 8'he1 == _t_T_74[15:8] ? 8'hf8 : _GEN_9440; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9442 = 8'he2 == _t_T_74[15:8] ? 8'h98 : _GEN_9441; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9443 = 8'he3 == _t_T_74[15:8] ? 8'h11 : _GEN_9442; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9444 = 8'he4 == _t_T_74[15:8] ? 8'h69 : _GEN_9443; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9445 = 8'he5 == _t_T_74[15:8] ? 8'hd9 : _GEN_9444; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9446 = 8'he6 == _t_T_74[15:8] ? 8'h8e : _GEN_9445; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9447 = 8'he7 == _t_T_74[15:8] ? 8'h94 : _GEN_9446; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9448 = 8'he8 == _t_T_74[15:8] ? 8'h9b : _GEN_9447; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9449 = 8'he9 == _t_T_74[15:8] ? 8'h1e : _GEN_9448; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9450 = 8'hea == _t_T_74[15:8] ? 8'h87 : _GEN_9449; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9451 = 8'heb == _t_T_74[15:8] ? 8'he9 : _GEN_9450; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9452 = 8'hec == _t_T_74[15:8] ? 8'hce : _GEN_9451; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9453 = 8'hed == _t_T_74[15:8] ? 8'h55 : _GEN_9452; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9454 = 8'hee == _t_T_74[15:8] ? 8'h28 : _GEN_9453; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9455 = 8'hef == _t_T_74[15:8] ? 8'hdf : _GEN_9454; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9456 = 8'hf0 == _t_T_74[15:8] ? 8'h8c : _GEN_9455; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9457 = 8'hf1 == _t_T_74[15:8] ? 8'ha1 : _GEN_9456; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9458 = 8'hf2 == _t_T_74[15:8] ? 8'h89 : _GEN_9457; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9459 = 8'hf3 == _t_T_74[15:8] ? 8'hd : _GEN_9458; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9460 = 8'hf4 == _t_T_74[15:8] ? 8'hbf : _GEN_9459; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9461 = 8'hf5 == _t_T_74[15:8] ? 8'he6 : _GEN_9460; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9462 = 8'hf6 == _t_T_74[15:8] ? 8'h42 : _GEN_9461; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9463 = 8'hf7 == _t_T_74[15:8] ? 8'h68 : _GEN_9462; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9464 = 8'hf8 == _t_T_74[15:8] ? 8'h41 : _GEN_9463; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9465 = 8'hf9 == _t_T_74[15:8] ? 8'h99 : _GEN_9464; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9466 = 8'hfa == _t_T_74[15:8] ? 8'h2d : _GEN_9465; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9467 = 8'hfb == _t_T_74[15:8] ? 8'hf : _GEN_9466; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9468 = 8'hfc == _t_T_74[15:8] ? 8'hb0 : _GEN_9467; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9469 = 8'hfd == _t_T_74[15:8] ? 8'h54 : _GEN_9468; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9470 = 8'hfe == _t_T_74[15:8] ? 8'hbb : _GEN_9469; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9471 = 8'hff == _t_T_74[15:8] ? 8'h16 : _GEN_9470; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9473 = 8'h1 == _t_T_74[7:0] ? 8'h7c : 8'h63; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9474 = 8'h2 == _t_T_74[7:0] ? 8'h77 : _GEN_9473; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9475 = 8'h3 == _t_T_74[7:0] ? 8'h7b : _GEN_9474; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9476 = 8'h4 == _t_T_74[7:0] ? 8'hf2 : _GEN_9475; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9477 = 8'h5 == _t_T_74[7:0] ? 8'h6b : _GEN_9476; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9478 = 8'h6 == _t_T_74[7:0] ? 8'h6f : _GEN_9477; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9479 = 8'h7 == _t_T_74[7:0] ? 8'hc5 : _GEN_9478; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9480 = 8'h8 == _t_T_74[7:0] ? 8'h30 : _GEN_9479; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9481 = 8'h9 == _t_T_74[7:0] ? 8'h1 : _GEN_9480; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9482 = 8'ha == _t_T_74[7:0] ? 8'h67 : _GEN_9481; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9483 = 8'hb == _t_T_74[7:0] ? 8'h2b : _GEN_9482; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9484 = 8'hc == _t_T_74[7:0] ? 8'hfe : _GEN_9483; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9485 = 8'hd == _t_T_74[7:0] ? 8'hd7 : _GEN_9484; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9486 = 8'he == _t_T_74[7:0] ? 8'hab : _GEN_9485; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9487 = 8'hf == _t_T_74[7:0] ? 8'h76 : _GEN_9486; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9488 = 8'h10 == _t_T_74[7:0] ? 8'hca : _GEN_9487; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9489 = 8'h11 == _t_T_74[7:0] ? 8'h82 : _GEN_9488; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9490 = 8'h12 == _t_T_74[7:0] ? 8'hc9 : _GEN_9489; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9491 = 8'h13 == _t_T_74[7:0] ? 8'h7d : _GEN_9490; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9492 = 8'h14 == _t_T_74[7:0] ? 8'hfa : _GEN_9491; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9493 = 8'h15 == _t_T_74[7:0] ? 8'h59 : _GEN_9492; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9494 = 8'h16 == _t_T_74[7:0] ? 8'h47 : _GEN_9493; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9495 = 8'h17 == _t_T_74[7:0] ? 8'hf0 : _GEN_9494; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9496 = 8'h18 == _t_T_74[7:0] ? 8'had : _GEN_9495; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9497 = 8'h19 == _t_T_74[7:0] ? 8'hd4 : _GEN_9496; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9498 = 8'h1a == _t_T_74[7:0] ? 8'ha2 : _GEN_9497; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9499 = 8'h1b == _t_T_74[7:0] ? 8'haf : _GEN_9498; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9500 = 8'h1c == _t_T_74[7:0] ? 8'h9c : _GEN_9499; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9501 = 8'h1d == _t_T_74[7:0] ? 8'ha4 : _GEN_9500; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9502 = 8'h1e == _t_T_74[7:0] ? 8'h72 : _GEN_9501; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9503 = 8'h1f == _t_T_74[7:0] ? 8'hc0 : _GEN_9502; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9504 = 8'h20 == _t_T_74[7:0] ? 8'hb7 : _GEN_9503; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9505 = 8'h21 == _t_T_74[7:0] ? 8'hfd : _GEN_9504; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9506 = 8'h22 == _t_T_74[7:0] ? 8'h93 : _GEN_9505; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9507 = 8'h23 == _t_T_74[7:0] ? 8'h26 : _GEN_9506; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9508 = 8'h24 == _t_T_74[7:0] ? 8'h36 : _GEN_9507; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9509 = 8'h25 == _t_T_74[7:0] ? 8'h3f : _GEN_9508; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9510 = 8'h26 == _t_T_74[7:0] ? 8'hf7 : _GEN_9509; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9511 = 8'h27 == _t_T_74[7:0] ? 8'hcc : _GEN_9510; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9512 = 8'h28 == _t_T_74[7:0] ? 8'h34 : _GEN_9511; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9513 = 8'h29 == _t_T_74[7:0] ? 8'ha5 : _GEN_9512; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9514 = 8'h2a == _t_T_74[7:0] ? 8'he5 : _GEN_9513; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9515 = 8'h2b == _t_T_74[7:0] ? 8'hf1 : _GEN_9514; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9516 = 8'h2c == _t_T_74[7:0] ? 8'h71 : _GEN_9515; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9517 = 8'h2d == _t_T_74[7:0] ? 8'hd8 : _GEN_9516; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9518 = 8'h2e == _t_T_74[7:0] ? 8'h31 : _GEN_9517; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9519 = 8'h2f == _t_T_74[7:0] ? 8'h15 : _GEN_9518; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9520 = 8'h30 == _t_T_74[7:0] ? 8'h4 : _GEN_9519; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9521 = 8'h31 == _t_T_74[7:0] ? 8'hc7 : _GEN_9520; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9522 = 8'h32 == _t_T_74[7:0] ? 8'h23 : _GEN_9521; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9523 = 8'h33 == _t_T_74[7:0] ? 8'hc3 : _GEN_9522; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9524 = 8'h34 == _t_T_74[7:0] ? 8'h18 : _GEN_9523; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9525 = 8'h35 == _t_T_74[7:0] ? 8'h96 : _GEN_9524; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9526 = 8'h36 == _t_T_74[7:0] ? 8'h5 : _GEN_9525; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9527 = 8'h37 == _t_T_74[7:0] ? 8'h9a : _GEN_9526; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9528 = 8'h38 == _t_T_74[7:0] ? 8'h7 : _GEN_9527; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9529 = 8'h39 == _t_T_74[7:0] ? 8'h12 : _GEN_9528; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9530 = 8'h3a == _t_T_74[7:0] ? 8'h80 : _GEN_9529; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9531 = 8'h3b == _t_T_74[7:0] ? 8'he2 : _GEN_9530; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9532 = 8'h3c == _t_T_74[7:0] ? 8'heb : _GEN_9531; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9533 = 8'h3d == _t_T_74[7:0] ? 8'h27 : _GEN_9532; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9534 = 8'h3e == _t_T_74[7:0] ? 8'hb2 : _GEN_9533; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9535 = 8'h3f == _t_T_74[7:0] ? 8'h75 : _GEN_9534; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9536 = 8'h40 == _t_T_74[7:0] ? 8'h9 : _GEN_9535; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9537 = 8'h41 == _t_T_74[7:0] ? 8'h83 : _GEN_9536; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9538 = 8'h42 == _t_T_74[7:0] ? 8'h2c : _GEN_9537; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9539 = 8'h43 == _t_T_74[7:0] ? 8'h1a : _GEN_9538; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9540 = 8'h44 == _t_T_74[7:0] ? 8'h1b : _GEN_9539; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9541 = 8'h45 == _t_T_74[7:0] ? 8'h6e : _GEN_9540; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9542 = 8'h46 == _t_T_74[7:0] ? 8'h5a : _GEN_9541; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9543 = 8'h47 == _t_T_74[7:0] ? 8'ha0 : _GEN_9542; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9544 = 8'h48 == _t_T_74[7:0] ? 8'h52 : _GEN_9543; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9545 = 8'h49 == _t_T_74[7:0] ? 8'h3b : _GEN_9544; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9546 = 8'h4a == _t_T_74[7:0] ? 8'hd6 : _GEN_9545; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9547 = 8'h4b == _t_T_74[7:0] ? 8'hb3 : _GEN_9546; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9548 = 8'h4c == _t_T_74[7:0] ? 8'h29 : _GEN_9547; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9549 = 8'h4d == _t_T_74[7:0] ? 8'he3 : _GEN_9548; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9550 = 8'h4e == _t_T_74[7:0] ? 8'h2f : _GEN_9549; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9551 = 8'h4f == _t_T_74[7:0] ? 8'h84 : _GEN_9550; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9552 = 8'h50 == _t_T_74[7:0] ? 8'h53 : _GEN_9551; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9553 = 8'h51 == _t_T_74[7:0] ? 8'hd1 : _GEN_9552; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9554 = 8'h52 == _t_T_74[7:0] ? 8'h0 : _GEN_9553; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9555 = 8'h53 == _t_T_74[7:0] ? 8'hed : _GEN_9554; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9556 = 8'h54 == _t_T_74[7:0] ? 8'h20 : _GEN_9555; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9557 = 8'h55 == _t_T_74[7:0] ? 8'hfc : _GEN_9556; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9558 = 8'h56 == _t_T_74[7:0] ? 8'hb1 : _GEN_9557; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9559 = 8'h57 == _t_T_74[7:0] ? 8'h5b : _GEN_9558; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9560 = 8'h58 == _t_T_74[7:0] ? 8'h6a : _GEN_9559; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9561 = 8'h59 == _t_T_74[7:0] ? 8'hcb : _GEN_9560; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9562 = 8'h5a == _t_T_74[7:0] ? 8'hbe : _GEN_9561; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9563 = 8'h5b == _t_T_74[7:0] ? 8'h39 : _GEN_9562; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9564 = 8'h5c == _t_T_74[7:0] ? 8'h4a : _GEN_9563; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9565 = 8'h5d == _t_T_74[7:0] ? 8'h4c : _GEN_9564; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9566 = 8'h5e == _t_T_74[7:0] ? 8'h58 : _GEN_9565; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9567 = 8'h5f == _t_T_74[7:0] ? 8'hcf : _GEN_9566; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9568 = 8'h60 == _t_T_74[7:0] ? 8'hd0 : _GEN_9567; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9569 = 8'h61 == _t_T_74[7:0] ? 8'hef : _GEN_9568; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9570 = 8'h62 == _t_T_74[7:0] ? 8'haa : _GEN_9569; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9571 = 8'h63 == _t_T_74[7:0] ? 8'hfb : _GEN_9570; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9572 = 8'h64 == _t_T_74[7:0] ? 8'h43 : _GEN_9571; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9573 = 8'h65 == _t_T_74[7:0] ? 8'h4d : _GEN_9572; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9574 = 8'h66 == _t_T_74[7:0] ? 8'h33 : _GEN_9573; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9575 = 8'h67 == _t_T_74[7:0] ? 8'h85 : _GEN_9574; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9576 = 8'h68 == _t_T_74[7:0] ? 8'h45 : _GEN_9575; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9577 = 8'h69 == _t_T_74[7:0] ? 8'hf9 : _GEN_9576; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9578 = 8'h6a == _t_T_74[7:0] ? 8'h2 : _GEN_9577; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9579 = 8'h6b == _t_T_74[7:0] ? 8'h7f : _GEN_9578; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9580 = 8'h6c == _t_T_74[7:0] ? 8'h50 : _GEN_9579; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9581 = 8'h6d == _t_T_74[7:0] ? 8'h3c : _GEN_9580; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9582 = 8'h6e == _t_T_74[7:0] ? 8'h9f : _GEN_9581; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9583 = 8'h6f == _t_T_74[7:0] ? 8'ha8 : _GEN_9582; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9584 = 8'h70 == _t_T_74[7:0] ? 8'h51 : _GEN_9583; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9585 = 8'h71 == _t_T_74[7:0] ? 8'ha3 : _GEN_9584; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9586 = 8'h72 == _t_T_74[7:0] ? 8'h40 : _GEN_9585; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9587 = 8'h73 == _t_T_74[7:0] ? 8'h8f : _GEN_9586; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9588 = 8'h74 == _t_T_74[7:0] ? 8'h92 : _GEN_9587; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9589 = 8'h75 == _t_T_74[7:0] ? 8'h9d : _GEN_9588; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9590 = 8'h76 == _t_T_74[7:0] ? 8'h38 : _GEN_9589; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9591 = 8'h77 == _t_T_74[7:0] ? 8'hf5 : _GEN_9590; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9592 = 8'h78 == _t_T_74[7:0] ? 8'hbc : _GEN_9591; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9593 = 8'h79 == _t_T_74[7:0] ? 8'hb6 : _GEN_9592; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9594 = 8'h7a == _t_T_74[7:0] ? 8'hda : _GEN_9593; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9595 = 8'h7b == _t_T_74[7:0] ? 8'h21 : _GEN_9594; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9596 = 8'h7c == _t_T_74[7:0] ? 8'h10 : _GEN_9595; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9597 = 8'h7d == _t_T_74[7:0] ? 8'hff : _GEN_9596; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9598 = 8'h7e == _t_T_74[7:0] ? 8'hf3 : _GEN_9597; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9599 = 8'h7f == _t_T_74[7:0] ? 8'hd2 : _GEN_9598; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9600 = 8'h80 == _t_T_74[7:0] ? 8'hcd : _GEN_9599; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9601 = 8'h81 == _t_T_74[7:0] ? 8'hc : _GEN_9600; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9602 = 8'h82 == _t_T_74[7:0] ? 8'h13 : _GEN_9601; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9603 = 8'h83 == _t_T_74[7:0] ? 8'hec : _GEN_9602; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9604 = 8'h84 == _t_T_74[7:0] ? 8'h5f : _GEN_9603; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9605 = 8'h85 == _t_T_74[7:0] ? 8'h97 : _GEN_9604; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9606 = 8'h86 == _t_T_74[7:0] ? 8'h44 : _GEN_9605; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9607 = 8'h87 == _t_T_74[7:0] ? 8'h17 : _GEN_9606; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9608 = 8'h88 == _t_T_74[7:0] ? 8'hc4 : _GEN_9607; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9609 = 8'h89 == _t_T_74[7:0] ? 8'ha7 : _GEN_9608; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9610 = 8'h8a == _t_T_74[7:0] ? 8'h7e : _GEN_9609; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9611 = 8'h8b == _t_T_74[7:0] ? 8'h3d : _GEN_9610; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9612 = 8'h8c == _t_T_74[7:0] ? 8'h64 : _GEN_9611; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9613 = 8'h8d == _t_T_74[7:0] ? 8'h5d : _GEN_9612; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9614 = 8'h8e == _t_T_74[7:0] ? 8'h19 : _GEN_9613; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9615 = 8'h8f == _t_T_74[7:0] ? 8'h73 : _GEN_9614; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9616 = 8'h90 == _t_T_74[7:0] ? 8'h60 : _GEN_9615; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9617 = 8'h91 == _t_T_74[7:0] ? 8'h81 : _GEN_9616; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9618 = 8'h92 == _t_T_74[7:0] ? 8'h4f : _GEN_9617; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9619 = 8'h93 == _t_T_74[7:0] ? 8'hdc : _GEN_9618; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9620 = 8'h94 == _t_T_74[7:0] ? 8'h22 : _GEN_9619; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9621 = 8'h95 == _t_T_74[7:0] ? 8'h2a : _GEN_9620; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9622 = 8'h96 == _t_T_74[7:0] ? 8'h90 : _GEN_9621; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9623 = 8'h97 == _t_T_74[7:0] ? 8'h88 : _GEN_9622; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9624 = 8'h98 == _t_T_74[7:0] ? 8'h46 : _GEN_9623; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9625 = 8'h99 == _t_T_74[7:0] ? 8'hee : _GEN_9624; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9626 = 8'h9a == _t_T_74[7:0] ? 8'hb8 : _GEN_9625; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9627 = 8'h9b == _t_T_74[7:0] ? 8'h14 : _GEN_9626; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9628 = 8'h9c == _t_T_74[7:0] ? 8'hde : _GEN_9627; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9629 = 8'h9d == _t_T_74[7:0] ? 8'h5e : _GEN_9628; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9630 = 8'h9e == _t_T_74[7:0] ? 8'hb : _GEN_9629; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9631 = 8'h9f == _t_T_74[7:0] ? 8'hdb : _GEN_9630; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9632 = 8'ha0 == _t_T_74[7:0] ? 8'he0 : _GEN_9631; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9633 = 8'ha1 == _t_T_74[7:0] ? 8'h32 : _GEN_9632; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9634 = 8'ha2 == _t_T_74[7:0] ? 8'h3a : _GEN_9633; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9635 = 8'ha3 == _t_T_74[7:0] ? 8'ha : _GEN_9634; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9636 = 8'ha4 == _t_T_74[7:0] ? 8'h49 : _GEN_9635; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9637 = 8'ha5 == _t_T_74[7:0] ? 8'h6 : _GEN_9636; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9638 = 8'ha6 == _t_T_74[7:0] ? 8'h24 : _GEN_9637; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9639 = 8'ha7 == _t_T_74[7:0] ? 8'h5c : _GEN_9638; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9640 = 8'ha8 == _t_T_74[7:0] ? 8'hc2 : _GEN_9639; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9641 = 8'ha9 == _t_T_74[7:0] ? 8'hd3 : _GEN_9640; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9642 = 8'haa == _t_T_74[7:0] ? 8'hac : _GEN_9641; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9643 = 8'hab == _t_T_74[7:0] ? 8'h62 : _GEN_9642; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9644 = 8'hac == _t_T_74[7:0] ? 8'h91 : _GEN_9643; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9645 = 8'had == _t_T_74[7:0] ? 8'h95 : _GEN_9644; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9646 = 8'hae == _t_T_74[7:0] ? 8'he4 : _GEN_9645; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9647 = 8'haf == _t_T_74[7:0] ? 8'h79 : _GEN_9646; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9648 = 8'hb0 == _t_T_74[7:0] ? 8'he7 : _GEN_9647; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9649 = 8'hb1 == _t_T_74[7:0] ? 8'hc8 : _GEN_9648; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9650 = 8'hb2 == _t_T_74[7:0] ? 8'h37 : _GEN_9649; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9651 = 8'hb3 == _t_T_74[7:0] ? 8'h6d : _GEN_9650; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9652 = 8'hb4 == _t_T_74[7:0] ? 8'h8d : _GEN_9651; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9653 = 8'hb5 == _t_T_74[7:0] ? 8'hd5 : _GEN_9652; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9654 = 8'hb6 == _t_T_74[7:0] ? 8'h4e : _GEN_9653; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9655 = 8'hb7 == _t_T_74[7:0] ? 8'ha9 : _GEN_9654; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9656 = 8'hb8 == _t_T_74[7:0] ? 8'h6c : _GEN_9655; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9657 = 8'hb9 == _t_T_74[7:0] ? 8'h56 : _GEN_9656; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9658 = 8'hba == _t_T_74[7:0] ? 8'hf4 : _GEN_9657; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9659 = 8'hbb == _t_T_74[7:0] ? 8'hea : _GEN_9658; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9660 = 8'hbc == _t_T_74[7:0] ? 8'h65 : _GEN_9659; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9661 = 8'hbd == _t_T_74[7:0] ? 8'h7a : _GEN_9660; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9662 = 8'hbe == _t_T_74[7:0] ? 8'hae : _GEN_9661; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9663 = 8'hbf == _t_T_74[7:0] ? 8'h8 : _GEN_9662; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9664 = 8'hc0 == _t_T_74[7:0] ? 8'hba : _GEN_9663; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9665 = 8'hc1 == _t_T_74[7:0] ? 8'h78 : _GEN_9664; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9666 = 8'hc2 == _t_T_74[7:0] ? 8'h25 : _GEN_9665; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9667 = 8'hc3 == _t_T_74[7:0] ? 8'h2e : _GEN_9666; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9668 = 8'hc4 == _t_T_74[7:0] ? 8'h1c : _GEN_9667; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9669 = 8'hc5 == _t_T_74[7:0] ? 8'ha6 : _GEN_9668; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9670 = 8'hc6 == _t_T_74[7:0] ? 8'hb4 : _GEN_9669; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9671 = 8'hc7 == _t_T_74[7:0] ? 8'hc6 : _GEN_9670; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9672 = 8'hc8 == _t_T_74[7:0] ? 8'he8 : _GEN_9671; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9673 = 8'hc9 == _t_T_74[7:0] ? 8'hdd : _GEN_9672; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9674 = 8'hca == _t_T_74[7:0] ? 8'h74 : _GEN_9673; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9675 = 8'hcb == _t_T_74[7:0] ? 8'h1f : _GEN_9674; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9676 = 8'hcc == _t_T_74[7:0] ? 8'h4b : _GEN_9675; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9677 = 8'hcd == _t_T_74[7:0] ? 8'hbd : _GEN_9676; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9678 = 8'hce == _t_T_74[7:0] ? 8'h8b : _GEN_9677; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9679 = 8'hcf == _t_T_74[7:0] ? 8'h8a : _GEN_9678; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9680 = 8'hd0 == _t_T_74[7:0] ? 8'h70 : _GEN_9679; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9681 = 8'hd1 == _t_T_74[7:0] ? 8'h3e : _GEN_9680; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9682 = 8'hd2 == _t_T_74[7:0] ? 8'hb5 : _GEN_9681; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9683 = 8'hd3 == _t_T_74[7:0] ? 8'h66 : _GEN_9682; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9684 = 8'hd4 == _t_T_74[7:0] ? 8'h48 : _GEN_9683; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9685 = 8'hd5 == _t_T_74[7:0] ? 8'h3 : _GEN_9684; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9686 = 8'hd6 == _t_T_74[7:0] ? 8'hf6 : _GEN_9685; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9687 = 8'hd7 == _t_T_74[7:0] ? 8'he : _GEN_9686; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9688 = 8'hd8 == _t_T_74[7:0] ? 8'h61 : _GEN_9687; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9689 = 8'hd9 == _t_T_74[7:0] ? 8'h35 : _GEN_9688; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9690 = 8'hda == _t_T_74[7:0] ? 8'h57 : _GEN_9689; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9691 = 8'hdb == _t_T_74[7:0] ? 8'hb9 : _GEN_9690; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9692 = 8'hdc == _t_T_74[7:0] ? 8'h86 : _GEN_9691; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9693 = 8'hdd == _t_T_74[7:0] ? 8'hc1 : _GEN_9692; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9694 = 8'hde == _t_T_74[7:0] ? 8'h1d : _GEN_9693; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9695 = 8'hdf == _t_T_74[7:0] ? 8'h9e : _GEN_9694; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9696 = 8'he0 == _t_T_74[7:0] ? 8'he1 : _GEN_9695; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9697 = 8'he1 == _t_T_74[7:0] ? 8'hf8 : _GEN_9696; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9698 = 8'he2 == _t_T_74[7:0] ? 8'h98 : _GEN_9697; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9699 = 8'he3 == _t_T_74[7:0] ? 8'h11 : _GEN_9698; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9700 = 8'he4 == _t_T_74[7:0] ? 8'h69 : _GEN_9699; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9701 = 8'he5 == _t_T_74[7:0] ? 8'hd9 : _GEN_9700; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9702 = 8'he6 == _t_T_74[7:0] ? 8'h8e : _GEN_9701; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9703 = 8'he7 == _t_T_74[7:0] ? 8'h94 : _GEN_9702; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9704 = 8'he8 == _t_T_74[7:0] ? 8'h9b : _GEN_9703; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9705 = 8'he9 == _t_T_74[7:0] ? 8'h1e : _GEN_9704; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9706 = 8'hea == _t_T_74[7:0] ? 8'h87 : _GEN_9705; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9707 = 8'heb == _t_T_74[7:0] ? 8'he9 : _GEN_9706; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9708 = 8'hec == _t_T_74[7:0] ? 8'hce : _GEN_9707; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9709 = 8'hed == _t_T_74[7:0] ? 8'h55 : _GEN_9708; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9710 = 8'hee == _t_T_74[7:0] ? 8'h28 : _GEN_9709; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9711 = 8'hef == _t_T_74[7:0] ? 8'hdf : _GEN_9710; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9712 = 8'hf0 == _t_T_74[7:0] ? 8'h8c : _GEN_9711; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9713 = 8'hf1 == _t_T_74[7:0] ? 8'ha1 : _GEN_9712; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9714 = 8'hf2 == _t_T_74[7:0] ? 8'h89 : _GEN_9713; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9715 = 8'hf3 == _t_T_74[7:0] ? 8'hd : _GEN_9714; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9716 = 8'hf4 == _t_T_74[7:0] ? 8'hbf : _GEN_9715; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9717 = 8'hf5 == _t_T_74[7:0] ? 8'he6 : _GEN_9716; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9718 = 8'hf6 == _t_T_74[7:0] ? 8'h42 : _GEN_9717; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9719 = 8'hf7 == _t_T_74[7:0] ? 8'h68 : _GEN_9718; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9720 = 8'hf8 == _t_T_74[7:0] ? 8'h41 : _GEN_9719; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9721 = 8'hf9 == _t_T_74[7:0] ? 8'h99 : _GEN_9720; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9722 = 8'hfa == _t_T_74[7:0] ? 8'h2d : _GEN_9721; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9723 = 8'hfb == _t_T_74[7:0] ? 8'hf : _GEN_9722; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9724 = 8'hfc == _t_T_74[7:0] ? 8'hb0 : _GEN_9723; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9725 = 8'hfd == _t_T_74[7:0] ? 8'h54 : _GEN_9724; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9726 = 8'hfe == _t_T_74[7:0] ? 8'hbb : _GEN_9725; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9727 = 8'hff == _t_T_74[7:0] ? 8'h16 : _GEN_9726; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9729 = 8'h1 == _t_T_74[31:24] ? 8'h7c : 8'h63; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9730 = 8'h2 == _t_T_74[31:24] ? 8'h77 : _GEN_9729; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9731 = 8'h3 == _t_T_74[31:24] ? 8'h7b : _GEN_9730; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9732 = 8'h4 == _t_T_74[31:24] ? 8'hf2 : _GEN_9731; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9733 = 8'h5 == _t_T_74[31:24] ? 8'h6b : _GEN_9732; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9734 = 8'h6 == _t_T_74[31:24] ? 8'h6f : _GEN_9733; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9735 = 8'h7 == _t_T_74[31:24] ? 8'hc5 : _GEN_9734; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9736 = 8'h8 == _t_T_74[31:24] ? 8'h30 : _GEN_9735; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9737 = 8'h9 == _t_T_74[31:24] ? 8'h1 : _GEN_9736; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9738 = 8'ha == _t_T_74[31:24] ? 8'h67 : _GEN_9737; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9739 = 8'hb == _t_T_74[31:24] ? 8'h2b : _GEN_9738; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9740 = 8'hc == _t_T_74[31:24] ? 8'hfe : _GEN_9739; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9741 = 8'hd == _t_T_74[31:24] ? 8'hd7 : _GEN_9740; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9742 = 8'he == _t_T_74[31:24] ? 8'hab : _GEN_9741; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9743 = 8'hf == _t_T_74[31:24] ? 8'h76 : _GEN_9742; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9744 = 8'h10 == _t_T_74[31:24] ? 8'hca : _GEN_9743; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9745 = 8'h11 == _t_T_74[31:24] ? 8'h82 : _GEN_9744; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9746 = 8'h12 == _t_T_74[31:24] ? 8'hc9 : _GEN_9745; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9747 = 8'h13 == _t_T_74[31:24] ? 8'h7d : _GEN_9746; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9748 = 8'h14 == _t_T_74[31:24] ? 8'hfa : _GEN_9747; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9749 = 8'h15 == _t_T_74[31:24] ? 8'h59 : _GEN_9748; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9750 = 8'h16 == _t_T_74[31:24] ? 8'h47 : _GEN_9749; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9751 = 8'h17 == _t_T_74[31:24] ? 8'hf0 : _GEN_9750; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9752 = 8'h18 == _t_T_74[31:24] ? 8'had : _GEN_9751; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9753 = 8'h19 == _t_T_74[31:24] ? 8'hd4 : _GEN_9752; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9754 = 8'h1a == _t_T_74[31:24] ? 8'ha2 : _GEN_9753; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9755 = 8'h1b == _t_T_74[31:24] ? 8'haf : _GEN_9754; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9756 = 8'h1c == _t_T_74[31:24] ? 8'h9c : _GEN_9755; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9757 = 8'h1d == _t_T_74[31:24] ? 8'ha4 : _GEN_9756; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9758 = 8'h1e == _t_T_74[31:24] ? 8'h72 : _GEN_9757; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9759 = 8'h1f == _t_T_74[31:24] ? 8'hc0 : _GEN_9758; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9760 = 8'h20 == _t_T_74[31:24] ? 8'hb7 : _GEN_9759; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9761 = 8'h21 == _t_T_74[31:24] ? 8'hfd : _GEN_9760; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9762 = 8'h22 == _t_T_74[31:24] ? 8'h93 : _GEN_9761; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9763 = 8'h23 == _t_T_74[31:24] ? 8'h26 : _GEN_9762; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9764 = 8'h24 == _t_T_74[31:24] ? 8'h36 : _GEN_9763; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9765 = 8'h25 == _t_T_74[31:24] ? 8'h3f : _GEN_9764; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9766 = 8'h26 == _t_T_74[31:24] ? 8'hf7 : _GEN_9765; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9767 = 8'h27 == _t_T_74[31:24] ? 8'hcc : _GEN_9766; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9768 = 8'h28 == _t_T_74[31:24] ? 8'h34 : _GEN_9767; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9769 = 8'h29 == _t_T_74[31:24] ? 8'ha5 : _GEN_9768; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9770 = 8'h2a == _t_T_74[31:24] ? 8'he5 : _GEN_9769; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9771 = 8'h2b == _t_T_74[31:24] ? 8'hf1 : _GEN_9770; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9772 = 8'h2c == _t_T_74[31:24] ? 8'h71 : _GEN_9771; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9773 = 8'h2d == _t_T_74[31:24] ? 8'hd8 : _GEN_9772; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9774 = 8'h2e == _t_T_74[31:24] ? 8'h31 : _GEN_9773; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9775 = 8'h2f == _t_T_74[31:24] ? 8'h15 : _GEN_9774; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9776 = 8'h30 == _t_T_74[31:24] ? 8'h4 : _GEN_9775; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9777 = 8'h31 == _t_T_74[31:24] ? 8'hc7 : _GEN_9776; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9778 = 8'h32 == _t_T_74[31:24] ? 8'h23 : _GEN_9777; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9779 = 8'h33 == _t_T_74[31:24] ? 8'hc3 : _GEN_9778; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9780 = 8'h34 == _t_T_74[31:24] ? 8'h18 : _GEN_9779; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9781 = 8'h35 == _t_T_74[31:24] ? 8'h96 : _GEN_9780; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9782 = 8'h36 == _t_T_74[31:24] ? 8'h5 : _GEN_9781; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9783 = 8'h37 == _t_T_74[31:24] ? 8'h9a : _GEN_9782; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9784 = 8'h38 == _t_T_74[31:24] ? 8'h7 : _GEN_9783; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9785 = 8'h39 == _t_T_74[31:24] ? 8'h12 : _GEN_9784; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9786 = 8'h3a == _t_T_74[31:24] ? 8'h80 : _GEN_9785; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9787 = 8'h3b == _t_T_74[31:24] ? 8'he2 : _GEN_9786; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9788 = 8'h3c == _t_T_74[31:24] ? 8'heb : _GEN_9787; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9789 = 8'h3d == _t_T_74[31:24] ? 8'h27 : _GEN_9788; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9790 = 8'h3e == _t_T_74[31:24] ? 8'hb2 : _GEN_9789; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9791 = 8'h3f == _t_T_74[31:24] ? 8'h75 : _GEN_9790; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9792 = 8'h40 == _t_T_74[31:24] ? 8'h9 : _GEN_9791; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9793 = 8'h41 == _t_T_74[31:24] ? 8'h83 : _GEN_9792; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9794 = 8'h42 == _t_T_74[31:24] ? 8'h2c : _GEN_9793; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9795 = 8'h43 == _t_T_74[31:24] ? 8'h1a : _GEN_9794; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9796 = 8'h44 == _t_T_74[31:24] ? 8'h1b : _GEN_9795; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9797 = 8'h45 == _t_T_74[31:24] ? 8'h6e : _GEN_9796; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9798 = 8'h46 == _t_T_74[31:24] ? 8'h5a : _GEN_9797; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9799 = 8'h47 == _t_T_74[31:24] ? 8'ha0 : _GEN_9798; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9800 = 8'h48 == _t_T_74[31:24] ? 8'h52 : _GEN_9799; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9801 = 8'h49 == _t_T_74[31:24] ? 8'h3b : _GEN_9800; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9802 = 8'h4a == _t_T_74[31:24] ? 8'hd6 : _GEN_9801; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9803 = 8'h4b == _t_T_74[31:24] ? 8'hb3 : _GEN_9802; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9804 = 8'h4c == _t_T_74[31:24] ? 8'h29 : _GEN_9803; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9805 = 8'h4d == _t_T_74[31:24] ? 8'he3 : _GEN_9804; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9806 = 8'h4e == _t_T_74[31:24] ? 8'h2f : _GEN_9805; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9807 = 8'h4f == _t_T_74[31:24] ? 8'h84 : _GEN_9806; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9808 = 8'h50 == _t_T_74[31:24] ? 8'h53 : _GEN_9807; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9809 = 8'h51 == _t_T_74[31:24] ? 8'hd1 : _GEN_9808; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9810 = 8'h52 == _t_T_74[31:24] ? 8'h0 : _GEN_9809; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9811 = 8'h53 == _t_T_74[31:24] ? 8'hed : _GEN_9810; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9812 = 8'h54 == _t_T_74[31:24] ? 8'h20 : _GEN_9811; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9813 = 8'h55 == _t_T_74[31:24] ? 8'hfc : _GEN_9812; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9814 = 8'h56 == _t_T_74[31:24] ? 8'hb1 : _GEN_9813; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9815 = 8'h57 == _t_T_74[31:24] ? 8'h5b : _GEN_9814; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9816 = 8'h58 == _t_T_74[31:24] ? 8'h6a : _GEN_9815; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9817 = 8'h59 == _t_T_74[31:24] ? 8'hcb : _GEN_9816; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9818 = 8'h5a == _t_T_74[31:24] ? 8'hbe : _GEN_9817; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9819 = 8'h5b == _t_T_74[31:24] ? 8'h39 : _GEN_9818; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9820 = 8'h5c == _t_T_74[31:24] ? 8'h4a : _GEN_9819; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9821 = 8'h5d == _t_T_74[31:24] ? 8'h4c : _GEN_9820; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9822 = 8'h5e == _t_T_74[31:24] ? 8'h58 : _GEN_9821; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9823 = 8'h5f == _t_T_74[31:24] ? 8'hcf : _GEN_9822; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9824 = 8'h60 == _t_T_74[31:24] ? 8'hd0 : _GEN_9823; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9825 = 8'h61 == _t_T_74[31:24] ? 8'hef : _GEN_9824; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9826 = 8'h62 == _t_T_74[31:24] ? 8'haa : _GEN_9825; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9827 = 8'h63 == _t_T_74[31:24] ? 8'hfb : _GEN_9826; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9828 = 8'h64 == _t_T_74[31:24] ? 8'h43 : _GEN_9827; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9829 = 8'h65 == _t_T_74[31:24] ? 8'h4d : _GEN_9828; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9830 = 8'h66 == _t_T_74[31:24] ? 8'h33 : _GEN_9829; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9831 = 8'h67 == _t_T_74[31:24] ? 8'h85 : _GEN_9830; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9832 = 8'h68 == _t_T_74[31:24] ? 8'h45 : _GEN_9831; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9833 = 8'h69 == _t_T_74[31:24] ? 8'hf9 : _GEN_9832; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9834 = 8'h6a == _t_T_74[31:24] ? 8'h2 : _GEN_9833; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9835 = 8'h6b == _t_T_74[31:24] ? 8'h7f : _GEN_9834; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9836 = 8'h6c == _t_T_74[31:24] ? 8'h50 : _GEN_9835; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9837 = 8'h6d == _t_T_74[31:24] ? 8'h3c : _GEN_9836; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9838 = 8'h6e == _t_T_74[31:24] ? 8'h9f : _GEN_9837; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9839 = 8'h6f == _t_T_74[31:24] ? 8'ha8 : _GEN_9838; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9840 = 8'h70 == _t_T_74[31:24] ? 8'h51 : _GEN_9839; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9841 = 8'h71 == _t_T_74[31:24] ? 8'ha3 : _GEN_9840; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9842 = 8'h72 == _t_T_74[31:24] ? 8'h40 : _GEN_9841; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9843 = 8'h73 == _t_T_74[31:24] ? 8'h8f : _GEN_9842; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9844 = 8'h74 == _t_T_74[31:24] ? 8'h92 : _GEN_9843; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9845 = 8'h75 == _t_T_74[31:24] ? 8'h9d : _GEN_9844; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9846 = 8'h76 == _t_T_74[31:24] ? 8'h38 : _GEN_9845; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9847 = 8'h77 == _t_T_74[31:24] ? 8'hf5 : _GEN_9846; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9848 = 8'h78 == _t_T_74[31:24] ? 8'hbc : _GEN_9847; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9849 = 8'h79 == _t_T_74[31:24] ? 8'hb6 : _GEN_9848; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9850 = 8'h7a == _t_T_74[31:24] ? 8'hda : _GEN_9849; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9851 = 8'h7b == _t_T_74[31:24] ? 8'h21 : _GEN_9850; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9852 = 8'h7c == _t_T_74[31:24] ? 8'h10 : _GEN_9851; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9853 = 8'h7d == _t_T_74[31:24] ? 8'hff : _GEN_9852; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9854 = 8'h7e == _t_T_74[31:24] ? 8'hf3 : _GEN_9853; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9855 = 8'h7f == _t_T_74[31:24] ? 8'hd2 : _GEN_9854; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9856 = 8'h80 == _t_T_74[31:24] ? 8'hcd : _GEN_9855; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9857 = 8'h81 == _t_T_74[31:24] ? 8'hc : _GEN_9856; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9858 = 8'h82 == _t_T_74[31:24] ? 8'h13 : _GEN_9857; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9859 = 8'h83 == _t_T_74[31:24] ? 8'hec : _GEN_9858; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9860 = 8'h84 == _t_T_74[31:24] ? 8'h5f : _GEN_9859; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9861 = 8'h85 == _t_T_74[31:24] ? 8'h97 : _GEN_9860; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9862 = 8'h86 == _t_T_74[31:24] ? 8'h44 : _GEN_9861; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9863 = 8'h87 == _t_T_74[31:24] ? 8'h17 : _GEN_9862; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9864 = 8'h88 == _t_T_74[31:24] ? 8'hc4 : _GEN_9863; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9865 = 8'h89 == _t_T_74[31:24] ? 8'ha7 : _GEN_9864; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9866 = 8'h8a == _t_T_74[31:24] ? 8'h7e : _GEN_9865; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9867 = 8'h8b == _t_T_74[31:24] ? 8'h3d : _GEN_9866; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9868 = 8'h8c == _t_T_74[31:24] ? 8'h64 : _GEN_9867; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9869 = 8'h8d == _t_T_74[31:24] ? 8'h5d : _GEN_9868; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9870 = 8'h8e == _t_T_74[31:24] ? 8'h19 : _GEN_9869; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9871 = 8'h8f == _t_T_74[31:24] ? 8'h73 : _GEN_9870; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9872 = 8'h90 == _t_T_74[31:24] ? 8'h60 : _GEN_9871; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9873 = 8'h91 == _t_T_74[31:24] ? 8'h81 : _GEN_9872; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9874 = 8'h92 == _t_T_74[31:24] ? 8'h4f : _GEN_9873; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9875 = 8'h93 == _t_T_74[31:24] ? 8'hdc : _GEN_9874; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9876 = 8'h94 == _t_T_74[31:24] ? 8'h22 : _GEN_9875; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9877 = 8'h95 == _t_T_74[31:24] ? 8'h2a : _GEN_9876; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9878 = 8'h96 == _t_T_74[31:24] ? 8'h90 : _GEN_9877; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9879 = 8'h97 == _t_T_74[31:24] ? 8'h88 : _GEN_9878; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9880 = 8'h98 == _t_T_74[31:24] ? 8'h46 : _GEN_9879; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9881 = 8'h99 == _t_T_74[31:24] ? 8'hee : _GEN_9880; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9882 = 8'h9a == _t_T_74[31:24] ? 8'hb8 : _GEN_9881; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9883 = 8'h9b == _t_T_74[31:24] ? 8'h14 : _GEN_9882; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9884 = 8'h9c == _t_T_74[31:24] ? 8'hde : _GEN_9883; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9885 = 8'h9d == _t_T_74[31:24] ? 8'h5e : _GEN_9884; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9886 = 8'h9e == _t_T_74[31:24] ? 8'hb : _GEN_9885; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9887 = 8'h9f == _t_T_74[31:24] ? 8'hdb : _GEN_9886; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9888 = 8'ha0 == _t_T_74[31:24] ? 8'he0 : _GEN_9887; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9889 = 8'ha1 == _t_T_74[31:24] ? 8'h32 : _GEN_9888; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9890 = 8'ha2 == _t_T_74[31:24] ? 8'h3a : _GEN_9889; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9891 = 8'ha3 == _t_T_74[31:24] ? 8'ha : _GEN_9890; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9892 = 8'ha4 == _t_T_74[31:24] ? 8'h49 : _GEN_9891; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9893 = 8'ha5 == _t_T_74[31:24] ? 8'h6 : _GEN_9892; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9894 = 8'ha6 == _t_T_74[31:24] ? 8'h24 : _GEN_9893; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9895 = 8'ha7 == _t_T_74[31:24] ? 8'h5c : _GEN_9894; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9896 = 8'ha8 == _t_T_74[31:24] ? 8'hc2 : _GEN_9895; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9897 = 8'ha9 == _t_T_74[31:24] ? 8'hd3 : _GEN_9896; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9898 = 8'haa == _t_T_74[31:24] ? 8'hac : _GEN_9897; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9899 = 8'hab == _t_T_74[31:24] ? 8'h62 : _GEN_9898; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9900 = 8'hac == _t_T_74[31:24] ? 8'h91 : _GEN_9899; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9901 = 8'had == _t_T_74[31:24] ? 8'h95 : _GEN_9900; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9902 = 8'hae == _t_T_74[31:24] ? 8'he4 : _GEN_9901; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9903 = 8'haf == _t_T_74[31:24] ? 8'h79 : _GEN_9902; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9904 = 8'hb0 == _t_T_74[31:24] ? 8'he7 : _GEN_9903; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9905 = 8'hb1 == _t_T_74[31:24] ? 8'hc8 : _GEN_9904; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9906 = 8'hb2 == _t_T_74[31:24] ? 8'h37 : _GEN_9905; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9907 = 8'hb3 == _t_T_74[31:24] ? 8'h6d : _GEN_9906; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9908 = 8'hb4 == _t_T_74[31:24] ? 8'h8d : _GEN_9907; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9909 = 8'hb5 == _t_T_74[31:24] ? 8'hd5 : _GEN_9908; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9910 = 8'hb6 == _t_T_74[31:24] ? 8'h4e : _GEN_9909; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9911 = 8'hb7 == _t_T_74[31:24] ? 8'ha9 : _GEN_9910; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9912 = 8'hb8 == _t_T_74[31:24] ? 8'h6c : _GEN_9911; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9913 = 8'hb9 == _t_T_74[31:24] ? 8'h56 : _GEN_9912; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9914 = 8'hba == _t_T_74[31:24] ? 8'hf4 : _GEN_9913; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9915 = 8'hbb == _t_T_74[31:24] ? 8'hea : _GEN_9914; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9916 = 8'hbc == _t_T_74[31:24] ? 8'h65 : _GEN_9915; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9917 = 8'hbd == _t_T_74[31:24] ? 8'h7a : _GEN_9916; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9918 = 8'hbe == _t_T_74[31:24] ? 8'hae : _GEN_9917; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9919 = 8'hbf == _t_T_74[31:24] ? 8'h8 : _GEN_9918; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9920 = 8'hc0 == _t_T_74[31:24] ? 8'hba : _GEN_9919; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9921 = 8'hc1 == _t_T_74[31:24] ? 8'h78 : _GEN_9920; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9922 = 8'hc2 == _t_T_74[31:24] ? 8'h25 : _GEN_9921; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9923 = 8'hc3 == _t_T_74[31:24] ? 8'h2e : _GEN_9922; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9924 = 8'hc4 == _t_T_74[31:24] ? 8'h1c : _GEN_9923; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9925 = 8'hc5 == _t_T_74[31:24] ? 8'ha6 : _GEN_9924; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9926 = 8'hc6 == _t_T_74[31:24] ? 8'hb4 : _GEN_9925; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9927 = 8'hc7 == _t_T_74[31:24] ? 8'hc6 : _GEN_9926; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9928 = 8'hc8 == _t_T_74[31:24] ? 8'he8 : _GEN_9927; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9929 = 8'hc9 == _t_T_74[31:24] ? 8'hdd : _GEN_9928; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9930 = 8'hca == _t_T_74[31:24] ? 8'h74 : _GEN_9929; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9931 = 8'hcb == _t_T_74[31:24] ? 8'h1f : _GEN_9930; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9932 = 8'hcc == _t_T_74[31:24] ? 8'h4b : _GEN_9931; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9933 = 8'hcd == _t_T_74[31:24] ? 8'hbd : _GEN_9932; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9934 = 8'hce == _t_T_74[31:24] ? 8'h8b : _GEN_9933; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9935 = 8'hcf == _t_T_74[31:24] ? 8'h8a : _GEN_9934; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9936 = 8'hd0 == _t_T_74[31:24] ? 8'h70 : _GEN_9935; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9937 = 8'hd1 == _t_T_74[31:24] ? 8'h3e : _GEN_9936; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9938 = 8'hd2 == _t_T_74[31:24] ? 8'hb5 : _GEN_9937; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9939 = 8'hd3 == _t_T_74[31:24] ? 8'h66 : _GEN_9938; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9940 = 8'hd4 == _t_T_74[31:24] ? 8'h48 : _GEN_9939; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9941 = 8'hd5 == _t_T_74[31:24] ? 8'h3 : _GEN_9940; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9942 = 8'hd6 == _t_T_74[31:24] ? 8'hf6 : _GEN_9941; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9943 = 8'hd7 == _t_T_74[31:24] ? 8'he : _GEN_9942; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9944 = 8'hd8 == _t_T_74[31:24] ? 8'h61 : _GEN_9943; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9945 = 8'hd9 == _t_T_74[31:24] ? 8'h35 : _GEN_9944; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9946 = 8'hda == _t_T_74[31:24] ? 8'h57 : _GEN_9945; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9947 = 8'hdb == _t_T_74[31:24] ? 8'hb9 : _GEN_9946; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9948 = 8'hdc == _t_T_74[31:24] ? 8'h86 : _GEN_9947; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9949 = 8'hdd == _t_T_74[31:24] ? 8'hc1 : _GEN_9948; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9950 = 8'hde == _t_T_74[31:24] ? 8'h1d : _GEN_9949; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9951 = 8'hdf == _t_T_74[31:24] ? 8'h9e : _GEN_9950; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9952 = 8'he0 == _t_T_74[31:24] ? 8'he1 : _GEN_9951; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9953 = 8'he1 == _t_T_74[31:24] ? 8'hf8 : _GEN_9952; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9954 = 8'he2 == _t_T_74[31:24] ? 8'h98 : _GEN_9953; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9955 = 8'he3 == _t_T_74[31:24] ? 8'h11 : _GEN_9954; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9956 = 8'he4 == _t_T_74[31:24] ? 8'h69 : _GEN_9955; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9957 = 8'he5 == _t_T_74[31:24] ? 8'hd9 : _GEN_9956; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9958 = 8'he6 == _t_T_74[31:24] ? 8'h8e : _GEN_9957; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9959 = 8'he7 == _t_T_74[31:24] ? 8'h94 : _GEN_9958; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9960 = 8'he8 == _t_T_74[31:24] ? 8'h9b : _GEN_9959; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9961 = 8'he9 == _t_T_74[31:24] ? 8'h1e : _GEN_9960; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9962 = 8'hea == _t_T_74[31:24] ? 8'h87 : _GEN_9961; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9963 = 8'heb == _t_T_74[31:24] ? 8'he9 : _GEN_9962; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9964 = 8'hec == _t_T_74[31:24] ? 8'hce : _GEN_9963; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9965 = 8'hed == _t_T_74[31:24] ? 8'h55 : _GEN_9964; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9966 = 8'hee == _t_T_74[31:24] ? 8'h28 : _GEN_9965; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9967 = 8'hef == _t_T_74[31:24] ? 8'hdf : _GEN_9966; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9968 = 8'hf0 == _t_T_74[31:24] ? 8'h8c : _GEN_9967; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9969 = 8'hf1 == _t_T_74[31:24] ? 8'ha1 : _GEN_9968; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9970 = 8'hf2 == _t_T_74[31:24] ? 8'h89 : _GEN_9969; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9971 = 8'hf3 == _t_T_74[31:24] ? 8'hd : _GEN_9970; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9972 = 8'hf4 == _t_T_74[31:24] ? 8'hbf : _GEN_9971; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9973 = 8'hf5 == _t_T_74[31:24] ? 8'he6 : _GEN_9972; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9974 = 8'hf6 == _t_T_74[31:24] ? 8'h42 : _GEN_9973; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9975 = 8'hf7 == _t_T_74[31:24] ? 8'h68 : _GEN_9974; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9976 = 8'hf8 == _t_T_74[31:24] ? 8'h41 : _GEN_9975; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9977 = 8'hf9 == _t_T_74[31:24] ? 8'h99 : _GEN_9976; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9978 = 8'hfa == _t_T_74[31:24] ? 8'h2d : _GEN_9977; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9979 = 8'hfb == _t_T_74[31:24] ? 8'hf : _GEN_9978; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9980 = 8'hfc == _t_T_74[31:24] ? 8'hb0 : _GEN_9979; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9981 = 8'hfd == _t_T_74[31:24] ? 8'h54 : _GEN_9980; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9982 = 8'hfe == _t_T_74[31:24] ? 8'hbb : _GEN_9981; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9983 = 8'hff == _t_T_74[31:24] ? 8'h16 : _GEN_9982; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9985 = 8'h1 == _t_T_74[23:16] ? 8'h7c : 8'h63; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9986 = 8'h2 == _t_T_74[23:16] ? 8'h77 : _GEN_9985; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9987 = 8'h3 == _t_T_74[23:16] ? 8'h7b : _GEN_9986; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9988 = 8'h4 == _t_T_74[23:16] ? 8'hf2 : _GEN_9987; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9989 = 8'h5 == _t_T_74[23:16] ? 8'h6b : _GEN_9988; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9990 = 8'h6 == _t_T_74[23:16] ? 8'h6f : _GEN_9989; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9991 = 8'h7 == _t_T_74[23:16] ? 8'hc5 : _GEN_9990; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9992 = 8'h8 == _t_T_74[23:16] ? 8'h30 : _GEN_9991; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9993 = 8'h9 == _t_T_74[23:16] ? 8'h1 : _GEN_9992; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9994 = 8'ha == _t_T_74[23:16] ? 8'h67 : _GEN_9993; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9995 = 8'hb == _t_T_74[23:16] ? 8'h2b : _GEN_9994; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9996 = 8'hc == _t_T_74[23:16] ? 8'hfe : _GEN_9995; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9997 = 8'hd == _t_T_74[23:16] ? 8'hd7 : _GEN_9996; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9998 = 8'he == _t_T_74[23:16] ? 8'hab : _GEN_9997; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_9999 = 8'hf == _t_T_74[23:16] ? 8'h76 : _GEN_9998; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10000 = 8'h10 == _t_T_74[23:16] ? 8'hca : _GEN_9999; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10001 = 8'h11 == _t_T_74[23:16] ? 8'h82 : _GEN_10000; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10002 = 8'h12 == _t_T_74[23:16] ? 8'hc9 : _GEN_10001; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10003 = 8'h13 == _t_T_74[23:16] ? 8'h7d : _GEN_10002; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10004 = 8'h14 == _t_T_74[23:16] ? 8'hfa : _GEN_10003; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10005 = 8'h15 == _t_T_74[23:16] ? 8'h59 : _GEN_10004; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10006 = 8'h16 == _t_T_74[23:16] ? 8'h47 : _GEN_10005; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10007 = 8'h17 == _t_T_74[23:16] ? 8'hf0 : _GEN_10006; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10008 = 8'h18 == _t_T_74[23:16] ? 8'had : _GEN_10007; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10009 = 8'h19 == _t_T_74[23:16] ? 8'hd4 : _GEN_10008; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10010 = 8'h1a == _t_T_74[23:16] ? 8'ha2 : _GEN_10009; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10011 = 8'h1b == _t_T_74[23:16] ? 8'haf : _GEN_10010; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10012 = 8'h1c == _t_T_74[23:16] ? 8'h9c : _GEN_10011; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10013 = 8'h1d == _t_T_74[23:16] ? 8'ha4 : _GEN_10012; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10014 = 8'h1e == _t_T_74[23:16] ? 8'h72 : _GEN_10013; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10015 = 8'h1f == _t_T_74[23:16] ? 8'hc0 : _GEN_10014; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10016 = 8'h20 == _t_T_74[23:16] ? 8'hb7 : _GEN_10015; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10017 = 8'h21 == _t_T_74[23:16] ? 8'hfd : _GEN_10016; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10018 = 8'h22 == _t_T_74[23:16] ? 8'h93 : _GEN_10017; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10019 = 8'h23 == _t_T_74[23:16] ? 8'h26 : _GEN_10018; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10020 = 8'h24 == _t_T_74[23:16] ? 8'h36 : _GEN_10019; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10021 = 8'h25 == _t_T_74[23:16] ? 8'h3f : _GEN_10020; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10022 = 8'h26 == _t_T_74[23:16] ? 8'hf7 : _GEN_10021; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10023 = 8'h27 == _t_T_74[23:16] ? 8'hcc : _GEN_10022; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10024 = 8'h28 == _t_T_74[23:16] ? 8'h34 : _GEN_10023; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10025 = 8'h29 == _t_T_74[23:16] ? 8'ha5 : _GEN_10024; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10026 = 8'h2a == _t_T_74[23:16] ? 8'he5 : _GEN_10025; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10027 = 8'h2b == _t_T_74[23:16] ? 8'hf1 : _GEN_10026; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10028 = 8'h2c == _t_T_74[23:16] ? 8'h71 : _GEN_10027; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10029 = 8'h2d == _t_T_74[23:16] ? 8'hd8 : _GEN_10028; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10030 = 8'h2e == _t_T_74[23:16] ? 8'h31 : _GEN_10029; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10031 = 8'h2f == _t_T_74[23:16] ? 8'h15 : _GEN_10030; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10032 = 8'h30 == _t_T_74[23:16] ? 8'h4 : _GEN_10031; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10033 = 8'h31 == _t_T_74[23:16] ? 8'hc7 : _GEN_10032; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10034 = 8'h32 == _t_T_74[23:16] ? 8'h23 : _GEN_10033; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10035 = 8'h33 == _t_T_74[23:16] ? 8'hc3 : _GEN_10034; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10036 = 8'h34 == _t_T_74[23:16] ? 8'h18 : _GEN_10035; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10037 = 8'h35 == _t_T_74[23:16] ? 8'h96 : _GEN_10036; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10038 = 8'h36 == _t_T_74[23:16] ? 8'h5 : _GEN_10037; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10039 = 8'h37 == _t_T_74[23:16] ? 8'h9a : _GEN_10038; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10040 = 8'h38 == _t_T_74[23:16] ? 8'h7 : _GEN_10039; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10041 = 8'h39 == _t_T_74[23:16] ? 8'h12 : _GEN_10040; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10042 = 8'h3a == _t_T_74[23:16] ? 8'h80 : _GEN_10041; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10043 = 8'h3b == _t_T_74[23:16] ? 8'he2 : _GEN_10042; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10044 = 8'h3c == _t_T_74[23:16] ? 8'heb : _GEN_10043; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10045 = 8'h3d == _t_T_74[23:16] ? 8'h27 : _GEN_10044; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10046 = 8'h3e == _t_T_74[23:16] ? 8'hb2 : _GEN_10045; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10047 = 8'h3f == _t_T_74[23:16] ? 8'h75 : _GEN_10046; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10048 = 8'h40 == _t_T_74[23:16] ? 8'h9 : _GEN_10047; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10049 = 8'h41 == _t_T_74[23:16] ? 8'h83 : _GEN_10048; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10050 = 8'h42 == _t_T_74[23:16] ? 8'h2c : _GEN_10049; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10051 = 8'h43 == _t_T_74[23:16] ? 8'h1a : _GEN_10050; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10052 = 8'h44 == _t_T_74[23:16] ? 8'h1b : _GEN_10051; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10053 = 8'h45 == _t_T_74[23:16] ? 8'h6e : _GEN_10052; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10054 = 8'h46 == _t_T_74[23:16] ? 8'h5a : _GEN_10053; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10055 = 8'h47 == _t_T_74[23:16] ? 8'ha0 : _GEN_10054; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10056 = 8'h48 == _t_T_74[23:16] ? 8'h52 : _GEN_10055; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10057 = 8'h49 == _t_T_74[23:16] ? 8'h3b : _GEN_10056; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10058 = 8'h4a == _t_T_74[23:16] ? 8'hd6 : _GEN_10057; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10059 = 8'h4b == _t_T_74[23:16] ? 8'hb3 : _GEN_10058; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10060 = 8'h4c == _t_T_74[23:16] ? 8'h29 : _GEN_10059; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10061 = 8'h4d == _t_T_74[23:16] ? 8'he3 : _GEN_10060; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10062 = 8'h4e == _t_T_74[23:16] ? 8'h2f : _GEN_10061; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10063 = 8'h4f == _t_T_74[23:16] ? 8'h84 : _GEN_10062; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10064 = 8'h50 == _t_T_74[23:16] ? 8'h53 : _GEN_10063; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10065 = 8'h51 == _t_T_74[23:16] ? 8'hd1 : _GEN_10064; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10066 = 8'h52 == _t_T_74[23:16] ? 8'h0 : _GEN_10065; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10067 = 8'h53 == _t_T_74[23:16] ? 8'hed : _GEN_10066; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10068 = 8'h54 == _t_T_74[23:16] ? 8'h20 : _GEN_10067; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10069 = 8'h55 == _t_T_74[23:16] ? 8'hfc : _GEN_10068; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10070 = 8'h56 == _t_T_74[23:16] ? 8'hb1 : _GEN_10069; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10071 = 8'h57 == _t_T_74[23:16] ? 8'h5b : _GEN_10070; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10072 = 8'h58 == _t_T_74[23:16] ? 8'h6a : _GEN_10071; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10073 = 8'h59 == _t_T_74[23:16] ? 8'hcb : _GEN_10072; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10074 = 8'h5a == _t_T_74[23:16] ? 8'hbe : _GEN_10073; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10075 = 8'h5b == _t_T_74[23:16] ? 8'h39 : _GEN_10074; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10076 = 8'h5c == _t_T_74[23:16] ? 8'h4a : _GEN_10075; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10077 = 8'h5d == _t_T_74[23:16] ? 8'h4c : _GEN_10076; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10078 = 8'h5e == _t_T_74[23:16] ? 8'h58 : _GEN_10077; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10079 = 8'h5f == _t_T_74[23:16] ? 8'hcf : _GEN_10078; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10080 = 8'h60 == _t_T_74[23:16] ? 8'hd0 : _GEN_10079; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10081 = 8'h61 == _t_T_74[23:16] ? 8'hef : _GEN_10080; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10082 = 8'h62 == _t_T_74[23:16] ? 8'haa : _GEN_10081; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10083 = 8'h63 == _t_T_74[23:16] ? 8'hfb : _GEN_10082; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10084 = 8'h64 == _t_T_74[23:16] ? 8'h43 : _GEN_10083; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10085 = 8'h65 == _t_T_74[23:16] ? 8'h4d : _GEN_10084; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10086 = 8'h66 == _t_T_74[23:16] ? 8'h33 : _GEN_10085; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10087 = 8'h67 == _t_T_74[23:16] ? 8'h85 : _GEN_10086; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10088 = 8'h68 == _t_T_74[23:16] ? 8'h45 : _GEN_10087; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10089 = 8'h69 == _t_T_74[23:16] ? 8'hf9 : _GEN_10088; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10090 = 8'h6a == _t_T_74[23:16] ? 8'h2 : _GEN_10089; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10091 = 8'h6b == _t_T_74[23:16] ? 8'h7f : _GEN_10090; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10092 = 8'h6c == _t_T_74[23:16] ? 8'h50 : _GEN_10091; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10093 = 8'h6d == _t_T_74[23:16] ? 8'h3c : _GEN_10092; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10094 = 8'h6e == _t_T_74[23:16] ? 8'h9f : _GEN_10093; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10095 = 8'h6f == _t_T_74[23:16] ? 8'ha8 : _GEN_10094; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10096 = 8'h70 == _t_T_74[23:16] ? 8'h51 : _GEN_10095; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10097 = 8'h71 == _t_T_74[23:16] ? 8'ha3 : _GEN_10096; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10098 = 8'h72 == _t_T_74[23:16] ? 8'h40 : _GEN_10097; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10099 = 8'h73 == _t_T_74[23:16] ? 8'h8f : _GEN_10098; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10100 = 8'h74 == _t_T_74[23:16] ? 8'h92 : _GEN_10099; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10101 = 8'h75 == _t_T_74[23:16] ? 8'h9d : _GEN_10100; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10102 = 8'h76 == _t_T_74[23:16] ? 8'h38 : _GEN_10101; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10103 = 8'h77 == _t_T_74[23:16] ? 8'hf5 : _GEN_10102; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10104 = 8'h78 == _t_T_74[23:16] ? 8'hbc : _GEN_10103; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10105 = 8'h79 == _t_T_74[23:16] ? 8'hb6 : _GEN_10104; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10106 = 8'h7a == _t_T_74[23:16] ? 8'hda : _GEN_10105; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10107 = 8'h7b == _t_T_74[23:16] ? 8'h21 : _GEN_10106; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10108 = 8'h7c == _t_T_74[23:16] ? 8'h10 : _GEN_10107; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10109 = 8'h7d == _t_T_74[23:16] ? 8'hff : _GEN_10108; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10110 = 8'h7e == _t_T_74[23:16] ? 8'hf3 : _GEN_10109; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10111 = 8'h7f == _t_T_74[23:16] ? 8'hd2 : _GEN_10110; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10112 = 8'h80 == _t_T_74[23:16] ? 8'hcd : _GEN_10111; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10113 = 8'h81 == _t_T_74[23:16] ? 8'hc : _GEN_10112; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10114 = 8'h82 == _t_T_74[23:16] ? 8'h13 : _GEN_10113; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10115 = 8'h83 == _t_T_74[23:16] ? 8'hec : _GEN_10114; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10116 = 8'h84 == _t_T_74[23:16] ? 8'h5f : _GEN_10115; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10117 = 8'h85 == _t_T_74[23:16] ? 8'h97 : _GEN_10116; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10118 = 8'h86 == _t_T_74[23:16] ? 8'h44 : _GEN_10117; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10119 = 8'h87 == _t_T_74[23:16] ? 8'h17 : _GEN_10118; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10120 = 8'h88 == _t_T_74[23:16] ? 8'hc4 : _GEN_10119; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10121 = 8'h89 == _t_T_74[23:16] ? 8'ha7 : _GEN_10120; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10122 = 8'h8a == _t_T_74[23:16] ? 8'h7e : _GEN_10121; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10123 = 8'h8b == _t_T_74[23:16] ? 8'h3d : _GEN_10122; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10124 = 8'h8c == _t_T_74[23:16] ? 8'h64 : _GEN_10123; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10125 = 8'h8d == _t_T_74[23:16] ? 8'h5d : _GEN_10124; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10126 = 8'h8e == _t_T_74[23:16] ? 8'h19 : _GEN_10125; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10127 = 8'h8f == _t_T_74[23:16] ? 8'h73 : _GEN_10126; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10128 = 8'h90 == _t_T_74[23:16] ? 8'h60 : _GEN_10127; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10129 = 8'h91 == _t_T_74[23:16] ? 8'h81 : _GEN_10128; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10130 = 8'h92 == _t_T_74[23:16] ? 8'h4f : _GEN_10129; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10131 = 8'h93 == _t_T_74[23:16] ? 8'hdc : _GEN_10130; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10132 = 8'h94 == _t_T_74[23:16] ? 8'h22 : _GEN_10131; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10133 = 8'h95 == _t_T_74[23:16] ? 8'h2a : _GEN_10132; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10134 = 8'h96 == _t_T_74[23:16] ? 8'h90 : _GEN_10133; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10135 = 8'h97 == _t_T_74[23:16] ? 8'h88 : _GEN_10134; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10136 = 8'h98 == _t_T_74[23:16] ? 8'h46 : _GEN_10135; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10137 = 8'h99 == _t_T_74[23:16] ? 8'hee : _GEN_10136; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10138 = 8'h9a == _t_T_74[23:16] ? 8'hb8 : _GEN_10137; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10139 = 8'h9b == _t_T_74[23:16] ? 8'h14 : _GEN_10138; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10140 = 8'h9c == _t_T_74[23:16] ? 8'hde : _GEN_10139; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10141 = 8'h9d == _t_T_74[23:16] ? 8'h5e : _GEN_10140; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10142 = 8'h9e == _t_T_74[23:16] ? 8'hb : _GEN_10141; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10143 = 8'h9f == _t_T_74[23:16] ? 8'hdb : _GEN_10142; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10144 = 8'ha0 == _t_T_74[23:16] ? 8'he0 : _GEN_10143; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10145 = 8'ha1 == _t_T_74[23:16] ? 8'h32 : _GEN_10144; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10146 = 8'ha2 == _t_T_74[23:16] ? 8'h3a : _GEN_10145; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10147 = 8'ha3 == _t_T_74[23:16] ? 8'ha : _GEN_10146; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10148 = 8'ha4 == _t_T_74[23:16] ? 8'h49 : _GEN_10147; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10149 = 8'ha5 == _t_T_74[23:16] ? 8'h6 : _GEN_10148; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10150 = 8'ha6 == _t_T_74[23:16] ? 8'h24 : _GEN_10149; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10151 = 8'ha7 == _t_T_74[23:16] ? 8'h5c : _GEN_10150; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10152 = 8'ha8 == _t_T_74[23:16] ? 8'hc2 : _GEN_10151; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10153 = 8'ha9 == _t_T_74[23:16] ? 8'hd3 : _GEN_10152; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10154 = 8'haa == _t_T_74[23:16] ? 8'hac : _GEN_10153; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10155 = 8'hab == _t_T_74[23:16] ? 8'h62 : _GEN_10154; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10156 = 8'hac == _t_T_74[23:16] ? 8'h91 : _GEN_10155; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10157 = 8'had == _t_T_74[23:16] ? 8'h95 : _GEN_10156; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10158 = 8'hae == _t_T_74[23:16] ? 8'he4 : _GEN_10157; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10159 = 8'haf == _t_T_74[23:16] ? 8'h79 : _GEN_10158; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10160 = 8'hb0 == _t_T_74[23:16] ? 8'he7 : _GEN_10159; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10161 = 8'hb1 == _t_T_74[23:16] ? 8'hc8 : _GEN_10160; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10162 = 8'hb2 == _t_T_74[23:16] ? 8'h37 : _GEN_10161; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10163 = 8'hb3 == _t_T_74[23:16] ? 8'h6d : _GEN_10162; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10164 = 8'hb4 == _t_T_74[23:16] ? 8'h8d : _GEN_10163; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10165 = 8'hb5 == _t_T_74[23:16] ? 8'hd5 : _GEN_10164; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10166 = 8'hb6 == _t_T_74[23:16] ? 8'h4e : _GEN_10165; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10167 = 8'hb7 == _t_T_74[23:16] ? 8'ha9 : _GEN_10166; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10168 = 8'hb8 == _t_T_74[23:16] ? 8'h6c : _GEN_10167; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10169 = 8'hb9 == _t_T_74[23:16] ? 8'h56 : _GEN_10168; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10170 = 8'hba == _t_T_74[23:16] ? 8'hf4 : _GEN_10169; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10171 = 8'hbb == _t_T_74[23:16] ? 8'hea : _GEN_10170; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10172 = 8'hbc == _t_T_74[23:16] ? 8'h65 : _GEN_10171; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10173 = 8'hbd == _t_T_74[23:16] ? 8'h7a : _GEN_10172; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10174 = 8'hbe == _t_T_74[23:16] ? 8'hae : _GEN_10173; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10175 = 8'hbf == _t_T_74[23:16] ? 8'h8 : _GEN_10174; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10176 = 8'hc0 == _t_T_74[23:16] ? 8'hba : _GEN_10175; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10177 = 8'hc1 == _t_T_74[23:16] ? 8'h78 : _GEN_10176; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10178 = 8'hc2 == _t_T_74[23:16] ? 8'h25 : _GEN_10177; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10179 = 8'hc3 == _t_T_74[23:16] ? 8'h2e : _GEN_10178; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10180 = 8'hc4 == _t_T_74[23:16] ? 8'h1c : _GEN_10179; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10181 = 8'hc5 == _t_T_74[23:16] ? 8'ha6 : _GEN_10180; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10182 = 8'hc6 == _t_T_74[23:16] ? 8'hb4 : _GEN_10181; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10183 = 8'hc7 == _t_T_74[23:16] ? 8'hc6 : _GEN_10182; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10184 = 8'hc8 == _t_T_74[23:16] ? 8'he8 : _GEN_10183; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10185 = 8'hc9 == _t_T_74[23:16] ? 8'hdd : _GEN_10184; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10186 = 8'hca == _t_T_74[23:16] ? 8'h74 : _GEN_10185; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10187 = 8'hcb == _t_T_74[23:16] ? 8'h1f : _GEN_10186; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10188 = 8'hcc == _t_T_74[23:16] ? 8'h4b : _GEN_10187; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10189 = 8'hcd == _t_T_74[23:16] ? 8'hbd : _GEN_10188; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10190 = 8'hce == _t_T_74[23:16] ? 8'h8b : _GEN_10189; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10191 = 8'hcf == _t_T_74[23:16] ? 8'h8a : _GEN_10190; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10192 = 8'hd0 == _t_T_74[23:16] ? 8'h70 : _GEN_10191; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10193 = 8'hd1 == _t_T_74[23:16] ? 8'h3e : _GEN_10192; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10194 = 8'hd2 == _t_T_74[23:16] ? 8'hb5 : _GEN_10193; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10195 = 8'hd3 == _t_T_74[23:16] ? 8'h66 : _GEN_10194; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10196 = 8'hd4 == _t_T_74[23:16] ? 8'h48 : _GEN_10195; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10197 = 8'hd5 == _t_T_74[23:16] ? 8'h3 : _GEN_10196; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10198 = 8'hd6 == _t_T_74[23:16] ? 8'hf6 : _GEN_10197; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10199 = 8'hd7 == _t_T_74[23:16] ? 8'he : _GEN_10198; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10200 = 8'hd8 == _t_T_74[23:16] ? 8'h61 : _GEN_10199; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10201 = 8'hd9 == _t_T_74[23:16] ? 8'h35 : _GEN_10200; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10202 = 8'hda == _t_T_74[23:16] ? 8'h57 : _GEN_10201; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10203 = 8'hdb == _t_T_74[23:16] ? 8'hb9 : _GEN_10202; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10204 = 8'hdc == _t_T_74[23:16] ? 8'h86 : _GEN_10203; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10205 = 8'hdd == _t_T_74[23:16] ? 8'hc1 : _GEN_10204; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10206 = 8'hde == _t_T_74[23:16] ? 8'h1d : _GEN_10205; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10207 = 8'hdf == _t_T_74[23:16] ? 8'h9e : _GEN_10206; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10208 = 8'he0 == _t_T_74[23:16] ? 8'he1 : _GEN_10207; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10209 = 8'he1 == _t_T_74[23:16] ? 8'hf8 : _GEN_10208; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10210 = 8'he2 == _t_T_74[23:16] ? 8'h98 : _GEN_10209; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10211 = 8'he3 == _t_T_74[23:16] ? 8'h11 : _GEN_10210; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10212 = 8'he4 == _t_T_74[23:16] ? 8'h69 : _GEN_10211; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10213 = 8'he5 == _t_T_74[23:16] ? 8'hd9 : _GEN_10212; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10214 = 8'he6 == _t_T_74[23:16] ? 8'h8e : _GEN_10213; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10215 = 8'he7 == _t_T_74[23:16] ? 8'h94 : _GEN_10214; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10216 = 8'he8 == _t_T_74[23:16] ? 8'h9b : _GEN_10215; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10217 = 8'he9 == _t_T_74[23:16] ? 8'h1e : _GEN_10216; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10218 = 8'hea == _t_T_74[23:16] ? 8'h87 : _GEN_10217; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10219 = 8'heb == _t_T_74[23:16] ? 8'he9 : _GEN_10218; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10220 = 8'hec == _t_T_74[23:16] ? 8'hce : _GEN_10219; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10221 = 8'hed == _t_T_74[23:16] ? 8'h55 : _GEN_10220; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10222 = 8'hee == _t_T_74[23:16] ? 8'h28 : _GEN_10221; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10223 = 8'hef == _t_T_74[23:16] ? 8'hdf : _GEN_10222; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10224 = 8'hf0 == _t_T_74[23:16] ? 8'h8c : _GEN_10223; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10225 = 8'hf1 == _t_T_74[23:16] ? 8'ha1 : _GEN_10224; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10226 = 8'hf2 == _t_T_74[23:16] ? 8'h89 : _GEN_10225; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10227 = 8'hf3 == _t_T_74[23:16] ? 8'hd : _GEN_10226; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10228 = 8'hf4 == _t_T_74[23:16] ? 8'hbf : _GEN_10227; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10229 = 8'hf5 == _t_T_74[23:16] ? 8'he6 : _GEN_10228; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10230 = 8'hf6 == _t_T_74[23:16] ? 8'h42 : _GEN_10229; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10231 = 8'hf7 == _t_T_74[23:16] ? 8'h68 : _GEN_10230; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10232 = 8'hf8 == _t_T_74[23:16] ? 8'h41 : _GEN_10231; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10233 = 8'hf9 == _t_T_74[23:16] ? 8'h99 : _GEN_10232; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10234 = 8'hfa == _t_T_74[23:16] ? 8'h2d : _GEN_10233; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10235 = 8'hfb == _t_T_74[23:16] ? 8'hf : _GEN_10234; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10236 = 8'hfc == _t_T_74[23:16] ? 8'hb0 : _GEN_10235; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10237 = 8'hfd == _t_T_74[23:16] ? 8'h54 : _GEN_10236; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10238 = 8'hfe == _t_T_74[23:16] ? 8'hbb : _GEN_10237; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [7:0] _GEN_10239 = 8'hff == _t_T_74[23:16] ? 8'h16 : _GEN_10238; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:{8,8}]
  wire [31:0] _t_T_79 = {_GEN_9983,_GEN_10239,_GEN_9471,_GEN_9727}; // @[src/main/scala/crypto/aes/KeySchedule.scala 26:8]
  wire [31:0] t_9 = _t_T_79 ^ 32'h36000000; // @[src/main/scala/crypto/aes/KeySchedule.scala 59:32]
  wire [31:0] w_40 = w_36 ^ t_9; // @[src/main/scala/crypto/aes/KeySchedule.scala 63:21]
  wire [31:0] w_41 = w_37 ^ w_40; // @[src/main/scala/crypto/aes/KeySchedule.scala 63:21]
  wire [31:0] w_42 = w_38 ^ w_41; // @[src/main/scala/crypto/aes/KeySchedule.scala 63:21]
  wire [31:0] w_43 = w_39 ^ w_42; // @[src/main/scala/crypto/aes/KeySchedule.scala 63:21]
  wire [63:0] io_rks_0_bits_lo = {w_2,w_3}; // @[src/main/scala/crypto/aes/KeySchedule.scala 75:26]
  wire [63:0] io_rks_0_bits_hi = {w_0,w_1}; // @[src/main/scala/crypto/aes/KeySchedule.scala 75:26]
  wire [63:0] io_rks_1_bits_lo = {w_6,w_7}; // @[src/main/scala/crypto/aes/KeySchedule.scala 75:26]
  wire [63:0] io_rks_1_bits_hi = {w_4,w_5}; // @[src/main/scala/crypto/aes/KeySchedule.scala 75:26]
  wire [63:0] io_rks_2_bits_lo = {w_10,w_11}; // @[src/main/scala/crypto/aes/KeySchedule.scala 75:26]
  wire [63:0] io_rks_2_bits_hi = {w_8,w_9}; // @[src/main/scala/crypto/aes/KeySchedule.scala 75:26]
  wire [63:0] io_rks_3_bits_lo = {w_14,w_15}; // @[src/main/scala/crypto/aes/KeySchedule.scala 75:26]
  wire [63:0] io_rks_3_bits_hi = {w_12,w_13}; // @[src/main/scala/crypto/aes/KeySchedule.scala 75:26]
  wire [63:0] io_rks_4_bits_lo = {w_18,w_19}; // @[src/main/scala/crypto/aes/KeySchedule.scala 75:26]
  wire [63:0] io_rks_4_bits_hi = {w_16,w_17}; // @[src/main/scala/crypto/aes/KeySchedule.scala 75:26]
  wire [63:0] io_rks_5_bits_lo = {w_22,w_23}; // @[src/main/scala/crypto/aes/KeySchedule.scala 75:26]
  wire [63:0] io_rks_5_bits_hi = {w_20,w_21}; // @[src/main/scala/crypto/aes/KeySchedule.scala 75:26]
  wire [63:0] io_rks_6_bits_lo = {w_26,w_27}; // @[src/main/scala/crypto/aes/KeySchedule.scala 75:26]
  wire [63:0] io_rks_6_bits_hi = {w_24,w_25}; // @[src/main/scala/crypto/aes/KeySchedule.scala 75:26]
  wire [63:0] io_rks_7_bits_lo = {w_30,w_31}; // @[src/main/scala/crypto/aes/KeySchedule.scala 75:26]
  wire [63:0] io_rks_7_bits_hi = {w_28,w_29}; // @[src/main/scala/crypto/aes/KeySchedule.scala 75:26]
  wire [63:0] io_rks_8_bits_lo = {w_34,w_35}; // @[src/main/scala/crypto/aes/KeySchedule.scala 75:26]
  wire [63:0] io_rks_8_bits_hi = {w_32,w_33}; // @[src/main/scala/crypto/aes/KeySchedule.scala 75:26]
  wire [63:0] io_rks_9_bits_lo = {w_38,w_39}; // @[src/main/scala/crypto/aes/KeySchedule.scala 75:26]
  wire [63:0] io_rks_9_bits_hi = {w_36,w_37}; // @[src/main/scala/crypto/aes/KeySchedule.scala 75:26]
  wire [63:0] io_rks_10_bits_lo = {w_42,w_43}; // @[src/main/scala/crypto/aes/KeySchedule.scala 75:26]
  wire [63:0] io_rks_10_bits_hi = {w_40,w_41}; // @[src/main/scala/crypto/aes/KeySchedule.scala 75:26]
  assign io_rks_0_bits = {io_rks_0_bits_hi,io_rks_0_bits_lo}; // @[src/main/scala/crypto/aes/KeySchedule.scala 75:26]
  assign io_rks_1_bits = {io_rks_1_bits_hi,io_rks_1_bits_lo}; // @[src/main/scala/crypto/aes/KeySchedule.scala 75:26]
  assign io_rks_2_bits = {io_rks_2_bits_hi,io_rks_2_bits_lo}; // @[src/main/scala/crypto/aes/KeySchedule.scala 75:26]
  assign io_rks_3_bits = {io_rks_3_bits_hi,io_rks_3_bits_lo}; // @[src/main/scala/crypto/aes/KeySchedule.scala 75:26]
  assign io_rks_4_bits = {io_rks_4_bits_hi,io_rks_4_bits_lo}; // @[src/main/scala/crypto/aes/KeySchedule.scala 75:26]
  assign io_rks_5_bits = {io_rks_5_bits_hi,io_rks_5_bits_lo}; // @[src/main/scala/crypto/aes/KeySchedule.scala 75:26]
  assign io_rks_6_bits = {io_rks_6_bits_hi,io_rks_6_bits_lo}; // @[src/main/scala/crypto/aes/KeySchedule.scala 75:26]
  assign io_rks_7_bits = {io_rks_7_bits_hi,io_rks_7_bits_lo}; // @[src/main/scala/crypto/aes/KeySchedule.scala 75:26]
  assign io_rks_8_bits = {io_rks_8_bits_hi,io_rks_8_bits_lo}; // @[src/main/scala/crypto/aes/KeySchedule.scala 75:26]
  assign io_rks_9_bits = {io_rks_9_bits_hi,io_rks_9_bits_lo}; // @[src/main/scala/crypto/aes/KeySchedule.scala 75:26]
  assign io_rks_10_bits = {io_rks_10_bits_hi,io_rks_10_bits_lo}; // @[src/main/scala/crypto/aes/KeySchedule.scala 75:26]
endmodule
module AddRoundKey(
  output         io_in_ready, // @[src/main/scala/crypto/aes/AddRoundKey.scala 21:29]
  input          io_in_valid, // @[src/main/scala/crypto/aes/AddRoundKey.scala 21:29]
  input  [127:0] io_in_bits_bits, // @[src/main/scala/crypto/aes/AddRoundKey.scala 21:29]
  input  [127:0] io_rk_bits, // @[src/main/scala/crypto/aes/AddRoundKey.scala 21:29]
  input          io_out_ready, // @[src/main/scala/crypto/aes/AddRoundKey.scala 21:29]
  output         io_out_valid, // @[src/main/scala/crypto/aes/AddRoundKey.scala 21:29]
  output [127:0] io_out_bits_bits // @[src/main/scala/crypto/aes/AddRoundKey.scala 21:29]
);
  assign io_in_ready = io_out_ready; // @[src/main/scala/crypto/aes/AddRoundKey.scala 25:16]
  assign io_out_valid = io_in_valid; // @[src/main/scala/crypto/aes/AddRoundKey.scala 24:16]
  assign io_out_bits_bits = io_in_bits_bits ^ io_rk_bits; // @[src/main/scala/crypto/aes/AddRoundKey.scala 26:39]
endmodule
module SubBytes(
  output         io_in_ready, // @[src/main/scala/crypto/aes/SubBytes.scala 9:14]
  input          io_in_valid, // @[src/main/scala/crypto/aes/SubBytes.scala 9:14]
  input  [127:0] io_in_bits_bits, // @[src/main/scala/crypto/aes/SubBytes.scala 9:14]
  input          io_out_ready, // @[src/main/scala/crypto/aes/SubBytes.scala 9:14]
  output         io_out_valid, // @[src/main/scala/crypto/aes/SubBytes.scala 9:14]
  output [127:0] io_out_bits_bits // @[src/main/scala/crypto/aes/SubBytes.scala 9:14]
);
  wire [7:0] inBytes_0 = io_in_bits_bits[127:120]; // @[src/main/scala/crypto/aes/SubBytes.scala 19:47]
  wire [7:0] inBytes_1 = io_in_bits_bits[119:112]; // @[src/main/scala/crypto/aes/SubBytes.scala 19:47]
  wire [7:0] inBytes_2 = io_in_bits_bits[111:104]; // @[src/main/scala/crypto/aes/SubBytes.scala 19:47]
  wire [7:0] inBytes_3 = io_in_bits_bits[103:96]; // @[src/main/scala/crypto/aes/SubBytes.scala 19:47]
  wire [7:0] inBytes_4 = io_in_bits_bits[95:88]; // @[src/main/scala/crypto/aes/SubBytes.scala 19:47]
  wire [7:0] inBytes_5 = io_in_bits_bits[87:80]; // @[src/main/scala/crypto/aes/SubBytes.scala 19:47]
  wire [7:0] inBytes_6 = io_in_bits_bits[79:72]; // @[src/main/scala/crypto/aes/SubBytes.scala 19:47]
  wire [7:0] inBytes_7 = io_in_bits_bits[71:64]; // @[src/main/scala/crypto/aes/SubBytes.scala 19:47]
  wire [7:0] inBytes_8 = io_in_bits_bits[63:56]; // @[src/main/scala/crypto/aes/SubBytes.scala 19:47]
  wire [7:0] inBytes_9 = io_in_bits_bits[55:48]; // @[src/main/scala/crypto/aes/SubBytes.scala 19:47]
  wire [7:0] inBytes_10 = io_in_bits_bits[47:40]; // @[src/main/scala/crypto/aes/SubBytes.scala 19:47]
  wire [7:0] inBytes_11 = io_in_bits_bits[39:32]; // @[src/main/scala/crypto/aes/SubBytes.scala 19:47]
  wire [7:0] inBytes_12 = io_in_bits_bits[31:24]; // @[src/main/scala/crypto/aes/SubBytes.scala 19:47]
  wire [7:0] inBytes_13 = io_in_bits_bits[23:16]; // @[src/main/scala/crypto/aes/SubBytes.scala 19:47]
  wire [7:0] inBytes_14 = io_in_bits_bits[15:8]; // @[src/main/scala/crypto/aes/SubBytes.scala 19:47]
  wire [7:0] inBytes_15 = io_in_bits_bits[7:0]; // @[src/main/scala/crypto/aes/SubBytes.scala 19:47]
  wire [7:0] _GEN_1 = 8'h1 == inBytes_0 ? 8'h7c : 8'h63; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2 = 8'h2 == inBytes_0 ? 8'h77 : _GEN_1; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3 = 8'h3 == inBytes_0 ? 8'h7b : _GEN_2; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_4 = 8'h4 == inBytes_0 ? 8'hf2 : _GEN_3; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_5 = 8'h5 == inBytes_0 ? 8'h6b : _GEN_4; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_6 = 8'h6 == inBytes_0 ? 8'h6f : _GEN_5; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_7 = 8'h7 == inBytes_0 ? 8'hc5 : _GEN_6; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_8 = 8'h8 == inBytes_0 ? 8'h30 : _GEN_7; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_9 = 8'h9 == inBytes_0 ? 8'h1 : _GEN_8; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_10 = 8'ha == inBytes_0 ? 8'h67 : _GEN_9; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_11 = 8'hb == inBytes_0 ? 8'h2b : _GEN_10; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_12 = 8'hc == inBytes_0 ? 8'hfe : _GEN_11; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_13 = 8'hd == inBytes_0 ? 8'hd7 : _GEN_12; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_14 = 8'he == inBytes_0 ? 8'hab : _GEN_13; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_15 = 8'hf == inBytes_0 ? 8'h76 : _GEN_14; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_16 = 8'h10 == inBytes_0 ? 8'hca : _GEN_15; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_17 = 8'h11 == inBytes_0 ? 8'h82 : _GEN_16; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_18 = 8'h12 == inBytes_0 ? 8'hc9 : _GEN_17; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_19 = 8'h13 == inBytes_0 ? 8'h7d : _GEN_18; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_20 = 8'h14 == inBytes_0 ? 8'hfa : _GEN_19; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_21 = 8'h15 == inBytes_0 ? 8'h59 : _GEN_20; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_22 = 8'h16 == inBytes_0 ? 8'h47 : _GEN_21; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_23 = 8'h17 == inBytes_0 ? 8'hf0 : _GEN_22; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_24 = 8'h18 == inBytes_0 ? 8'had : _GEN_23; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_25 = 8'h19 == inBytes_0 ? 8'hd4 : _GEN_24; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_26 = 8'h1a == inBytes_0 ? 8'ha2 : _GEN_25; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_27 = 8'h1b == inBytes_0 ? 8'haf : _GEN_26; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_28 = 8'h1c == inBytes_0 ? 8'h9c : _GEN_27; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_29 = 8'h1d == inBytes_0 ? 8'ha4 : _GEN_28; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_30 = 8'h1e == inBytes_0 ? 8'h72 : _GEN_29; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_31 = 8'h1f == inBytes_0 ? 8'hc0 : _GEN_30; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_32 = 8'h20 == inBytes_0 ? 8'hb7 : _GEN_31; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_33 = 8'h21 == inBytes_0 ? 8'hfd : _GEN_32; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_34 = 8'h22 == inBytes_0 ? 8'h93 : _GEN_33; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_35 = 8'h23 == inBytes_0 ? 8'h26 : _GEN_34; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_36 = 8'h24 == inBytes_0 ? 8'h36 : _GEN_35; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_37 = 8'h25 == inBytes_0 ? 8'h3f : _GEN_36; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_38 = 8'h26 == inBytes_0 ? 8'hf7 : _GEN_37; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_39 = 8'h27 == inBytes_0 ? 8'hcc : _GEN_38; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_40 = 8'h28 == inBytes_0 ? 8'h34 : _GEN_39; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_41 = 8'h29 == inBytes_0 ? 8'ha5 : _GEN_40; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_42 = 8'h2a == inBytes_0 ? 8'he5 : _GEN_41; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_43 = 8'h2b == inBytes_0 ? 8'hf1 : _GEN_42; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_44 = 8'h2c == inBytes_0 ? 8'h71 : _GEN_43; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_45 = 8'h2d == inBytes_0 ? 8'hd8 : _GEN_44; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_46 = 8'h2e == inBytes_0 ? 8'h31 : _GEN_45; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_47 = 8'h2f == inBytes_0 ? 8'h15 : _GEN_46; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_48 = 8'h30 == inBytes_0 ? 8'h4 : _GEN_47; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_49 = 8'h31 == inBytes_0 ? 8'hc7 : _GEN_48; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_50 = 8'h32 == inBytes_0 ? 8'h23 : _GEN_49; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_51 = 8'h33 == inBytes_0 ? 8'hc3 : _GEN_50; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_52 = 8'h34 == inBytes_0 ? 8'h18 : _GEN_51; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_53 = 8'h35 == inBytes_0 ? 8'h96 : _GEN_52; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_54 = 8'h36 == inBytes_0 ? 8'h5 : _GEN_53; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_55 = 8'h37 == inBytes_0 ? 8'h9a : _GEN_54; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_56 = 8'h38 == inBytes_0 ? 8'h7 : _GEN_55; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_57 = 8'h39 == inBytes_0 ? 8'h12 : _GEN_56; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_58 = 8'h3a == inBytes_0 ? 8'h80 : _GEN_57; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_59 = 8'h3b == inBytes_0 ? 8'he2 : _GEN_58; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_60 = 8'h3c == inBytes_0 ? 8'heb : _GEN_59; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_61 = 8'h3d == inBytes_0 ? 8'h27 : _GEN_60; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_62 = 8'h3e == inBytes_0 ? 8'hb2 : _GEN_61; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_63 = 8'h3f == inBytes_0 ? 8'h75 : _GEN_62; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_64 = 8'h40 == inBytes_0 ? 8'h9 : _GEN_63; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_65 = 8'h41 == inBytes_0 ? 8'h83 : _GEN_64; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_66 = 8'h42 == inBytes_0 ? 8'h2c : _GEN_65; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_67 = 8'h43 == inBytes_0 ? 8'h1a : _GEN_66; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_68 = 8'h44 == inBytes_0 ? 8'h1b : _GEN_67; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_69 = 8'h45 == inBytes_0 ? 8'h6e : _GEN_68; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_70 = 8'h46 == inBytes_0 ? 8'h5a : _GEN_69; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_71 = 8'h47 == inBytes_0 ? 8'ha0 : _GEN_70; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_72 = 8'h48 == inBytes_0 ? 8'h52 : _GEN_71; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_73 = 8'h49 == inBytes_0 ? 8'h3b : _GEN_72; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_74 = 8'h4a == inBytes_0 ? 8'hd6 : _GEN_73; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_75 = 8'h4b == inBytes_0 ? 8'hb3 : _GEN_74; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_76 = 8'h4c == inBytes_0 ? 8'h29 : _GEN_75; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_77 = 8'h4d == inBytes_0 ? 8'he3 : _GEN_76; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_78 = 8'h4e == inBytes_0 ? 8'h2f : _GEN_77; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_79 = 8'h4f == inBytes_0 ? 8'h84 : _GEN_78; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_80 = 8'h50 == inBytes_0 ? 8'h53 : _GEN_79; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_81 = 8'h51 == inBytes_0 ? 8'hd1 : _GEN_80; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_82 = 8'h52 == inBytes_0 ? 8'h0 : _GEN_81; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_83 = 8'h53 == inBytes_0 ? 8'hed : _GEN_82; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_84 = 8'h54 == inBytes_0 ? 8'h20 : _GEN_83; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_85 = 8'h55 == inBytes_0 ? 8'hfc : _GEN_84; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_86 = 8'h56 == inBytes_0 ? 8'hb1 : _GEN_85; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_87 = 8'h57 == inBytes_0 ? 8'h5b : _GEN_86; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_88 = 8'h58 == inBytes_0 ? 8'h6a : _GEN_87; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_89 = 8'h59 == inBytes_0 ? 8'hcb : _GEN_88; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_90 = 8'h5a == inBytes_0 ? 8'hbe : _GEN_89; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_91 = 8'h5b == inBytes_0 ? 8'h39 : _GEN_90; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_92 = 8'h5c == inBytes_0 ? 8'h4a : _GEN_91; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_93 = 8'h5d == inBytes_0 ? 8'h4c : _GEN_92; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_94 = 8'h5e == inBytes_0 ? 8'h58 : _GEN_93; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_95 = 8'h5f == inBytes_0 ? 8'hcf : _GEN_94; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_96 = 8'h60 == inBytes_0 ? 8'hd0 : _GEN_95; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_97 = 8'h61 == inBytes_0 ? 8'hef : _GEN_96; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_98 = 8'h62 == inBytes_0 ? 8'haa : _GEN_97; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_99 = 8'h63 == inBytes_0 ? 8'hfb : _GEN_98; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_100 = 8'h64 == inBytes_0 ? 8'h43 : _GEN_99; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_101 = 8'h65 == inBytes_0 ? 8'h4d : _GEN_100; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_102 = 8'h66 == inBytes_0 ? 8'h33 : _GEN_101; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_103 = 8'h67 == inBytes_0 ? 8'h85 : _GEN_102; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_104 = 8'h68 == inBytes_0 ? 8'h45 : _GEN_103; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_105 = 8'h69 == inBytes_0 ? 8'hf9 : _GEN_104; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_106 = 8'h6a == inBytes_0 ? 8'h2 : _GEN_105; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_107 = 8'h6b == inBytes_0 ? 8'h7f : _GEN_106; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_108 = 8'h6c == inBytes_0 ? 8'h50 : _GEN_107; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_109 = 8'h6d == inBytes_0 ? 8'h3c : _GEN_108; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_110 = 8'h6e == inBytes_0 ? 8'h9f : _GEN_109; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_111 = 8'h6f == inBytes_0 ? 8'ha8 : _GEN_110; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_112 = 8'h70 == inBytes_0 ? 8'h51 : _GEN_111; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_113 = 8'h71 == inBytes_0 ? 8'ha3 : _GEN_112; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_114 = 8'h72 == inBytes_0 ? 8'h40 : _GEN_113; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_115 = 8'h73 == inBytes_0 ? 8'h8f : _GEN_114; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_116 = 8'h74 == inBytes_0 ? 8'h92 : _GEN_115; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_117 = 8'h75 == inBytes_0 ? 8'h9d : _GEN_116; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_118 = 8'h76 == inBytes_0 ? 8'h38 : _GEN_117; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_119 = 8'h77 == inBytes_0 ? 8'hf5 : _GEN_118; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_120 = 8'h78 == inBytes_0 ? 8'hbc : _GEN_119; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_121 = 8'h79 == inBytes_0 ? 8'hb6 : _GEN_120; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_122 = 8'h7a == inBytes_0 ? 8'hda : _GEN_121; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_123 = 8'h7b == inBytes_0 ? 8'h21 : _GEN_122; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_124 = 8'h7c == inBytes_0 ? 8'h10 : _GEN_123; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_125 = 8'h7d == inBytes_0 ? 8'hff : _GEN_124; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_126 = 8'h7e == inBytes_0 ? 8'hf3 : _GEN_125; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_127 = 8'h7f == inBytes_0 ? 8'hd2 : _GEN_126; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_128 = 8'h80 == inBytes_0 ? 8'hcd : _GEN_127; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_129 = 8'h81 == inBytes_0 ? 8'hc : _GEN_128; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_130 = 8'h82 == inBytes_0 ? 8'h13 : _GEN_129; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_131 = 8'h83 == inBytes_0 ? 8'hec : _GEN_130; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_132 = 8'h84 == inBytes_0 ? 8'h5f : _GEN_131; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_133 = 8'h85 == inBytes_0 ? 8'h97 : _GEN_132; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_134 = 8'h86 == inBytes_0 ? 8'h44 : _GEN_133; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_135 = 8'h87 == inBytes_0 ? 8'h17 : _GEN_134; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_136 = 8'h88 == inBytes_0 ? 8'hc4 : _GEN_135; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_137 = 8'h89 == inBytes_0 ? 8'ha7 : _GEN_136; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_138 = 8'h8a == inBytes_0 ? 8'h7e : _GEN_137; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_139 = 8'h8b == inBytes_0 ? 8'h3d : _GEN_138; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_140 = 8'h8c == inBytes_0 ? 8'h64 : _GEN_139; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_141 = 8'h8d == inBytes_0 ? 8'h5d : _GEN_140; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_142 = 8'h8e == inBytes_0 ? 8'h19 : _GEN_141; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_143 = 8'h8f == inBytes_0 ? 8'h73 : _GEN_142; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_144 = 8'h90 == inBytes_0 ? 8'h60 : _GEN_143; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_145 = 8'h91 == inBytes_0 ? 8'h81 : _GEN_144; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_146 = 8'h92 == inBytes_0 ? 8'h4f : _GEN_145; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_147 = 8'h93 == inBytes_0 ? 8'hdc : _GEN_146; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_148 = 8'h94 == inBytes_0 ? 8'h22 : _GEN_147; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_149 = 8'h95 == inBytes_0 ? 8'h2a : _GEN_148; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_150 = 8'h96 == inBytes_0 ? 8'h90 : _GEN_149; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_151 = 8'h97 == inBytes_0 ? 8'h88 : _GEN_150; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_152 = 8'h98 == inBytes_0 ? 8'h46 : _GEN_151; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_153 = 8'h99 == inBytes_0 ? 8'hee : _GEN_152; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_154 = 8'h9a == inBytes_0 ? 8'hb8 : _GEN_153; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_155 = 8'h9b == inBytes_0 ? 8'h14 : _GEN_154; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_156 = 8'h9c == inBytes_0 ? 8'hde : _GEN_155; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_157 = 8'h9d == inBytes_0 ? 8'h5e : _GEN_156; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_158 = 8'h9e == inBytes_0 ? 8'hb : _GEN_157; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_159 = 8'h9f == inBytes_0 ? 8'hdb : _GEN_158; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_160 = 8'ha0 == inBytes_0 ? 8'he0 : _GEN_159; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_161 = 8'ha1 == inBytes_0 ? 8'h32 : _GEN_160; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_162 = 8'ha2 == inBytes_0 ? 8'h3a : _GEN_161; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_163 = 8'ha3 == inBytes_0 ? 8'ha : _GEN_162; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_164 = 8'ha4 == inBytes_0 ? 8'h49 : _GEN_163; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_165 = 8'ha5 == inBytes_0 ? 8'h6 : _GEN_164; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_166 = 8'ha6 == inBytes_0 ? 8'h24 : _GEN_165; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_167 = 8'ha7 == inBytes_0 ? 8'h5c : _GEN_166; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_168 = 8'ha8 == inBytes_0 ? 8'hc2 : _GEN_167; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_169 = 8'ha9 == inBytes_0 ? 8'hd3 : _GEN_168; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_170 = 8'haa == inBytes_0 ? 8'hac : _GEN_169; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_171 = 8'hab == inBytes_0 ? 8'h62 : _GEN_170; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_172 = 8'hac == inBytes_0 ? 8'h91 : _GEN_171; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_173 = 8'had == inBytes_0 ? 8'h95 : _GEN_172; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_174 = 8'hae == inBytes_0 ? 8'he4 : _GEN_173; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_175 = 8'haf == inBytes_0 ? 8'h79 : _GEN_174; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_176 = 8'hb0 == inBytes_0 ? 8'he7 : _GEN_175; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_177 = 8'hb1 == inBytes_0 ? 8'hc8 : _GEN_176; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_178 = 8'hb2 == inBytes_0 ? 8'h37 : _GEN_177; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_179 = 8'hb3 == inBytes_0 ? 8'h6d : _GEN_178; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_180 = 8'hb4 == inBytes_0 ? 8'h8d : _GEN_179; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_181 = 8'hb5 == inBytes_0 ? 8'hd5 : _GEN_180; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_182 = 8'hb6 == inBytes_0 ? 8'h4e : _GEN_181; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_183 = 8'hb7 == inBytes_0 ? 8'ha9 : _GEN_182; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_184 = 8'hb8 == inBytes_0 ? 8'h6c : _GEN_183; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_185 = 8'hb9 == inBytes_0 ? 8'h56 : _GEN_184; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_186 = 8'hba == inBytes_0 ? 8'hf4 : _GEN_185; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_187 = 8'hbb == inBytes_0 ? 8'hea : _GEN_186; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_188 = 8'hbc == inBytes_0 ? 8'h65 : _GEN_187; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_189 = 8'hbd == inBytes_0 ? 8'h7a : _GEN_188; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_190 = 8'hbe == inBytes_0 ? 8'hae : _GEN_189; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_191 = 8'hbf == inBytes_0 ? 8'h8 : _GEN_190; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_192 = 8'hc0 == inBytes_0 ? 8'hba : _GEN_191; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_193 = 8'hc1 == inBytes_0 ? 8'h78 : _GEN_192; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_194 = 8'hc2 == inBytes_0 ? 8'h25 : _GEN_193; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_195 = 8'hc3 == inBytes_0 ? 8'h2e : _GEN_194; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_196 = 8'hc4 == inBytes_0 ? 8'h1c : _GEN_195; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_197 = 8'hc5 == inBytes_0 ? 8'ha6 : _GEN_196; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_198 = 8'hc6 == inBytes_0 ? 8'hb4 : _GEN_197; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_199 = 8'hc7 == inBytes_0 ? 8'hc6 : _GEN_198; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_200 = 8'hc8 == inBytes_0 ? 8'he8 : _GEN_199; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_201 = 8'hc9 == inBytes_0 ? 8'hdd : _GEN_200; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_202 = 8'hca == inBytes_0 ? 8'h74 : _GEN_201; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_203 = 8'hcb == inBytes_0 ? 8'h1f : _GEN_202; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_204 = 8'hcc == inBytes_0 ? 8'h4b : _GEN_203; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_205 = 8'hcd == inBytes_0 ? 8'hbd : _GEN_204; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_206 = 8'hce == inBytes_0 ? 8'h8b : _GEN_205; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_207 = 8'hcf == inBytes_0 ? 8'h8a : _GEN_206; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_208 = 8'hd0 == inBytes_0 ? 8'h70 : _GEN_207; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_209 = 8'hd1 == inBytes_0 ? 8'h3e : _GEN_208; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_210 = 8'hd2 == inBytes_0 ? 8'hb5 : _GEN_209; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_211 = 8'hd3 == inBytes_0 ? 8'h66 : _GEN_210; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_212 = 8'hd4 == inBytes_0 ? 8'h48 : _GEN_211; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_213 = 8'hd5 == inBytes_0 ? 8'h3 : _GEN_212; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_214 = 8'hd6 == inBytes_0 ? 8'hf6 : _GEN_213; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_215 = 8'hd7 == inBytes_0 ? 8'he : _GEN_214; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_216 = 8'hd8 == inBytes_0 ? 8'h61 : _GEN_215; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_217 = 8'hd9 == inBytes_0 ? 8'h35 : _GEN_216; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_218 = 8'hda == inBytes_0 ? 8'h57 : _GEN_217; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_219 = 8'hdb == inBytes_0 ? 8'hb9 : _GEN_218; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_220 = 8'hdc == inBytes_0 ? 8'h86 : _GEN_219; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_221 = 8'hdd == inBytes_0 ? 8'hc1 : _GEN_220; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_222 = 8'hde == inBytes_0 ? 8'h1d : _GEN_221; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_223 = 8'hdf == inBytes_0 ? 8'h9e : _GEN_222; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_224 = 8'he0 == inBytes_0 ? 8'he1 : _GEN_223; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_225 = 8'he1 == inBytes_0 ? 8'hf8 : _GEN_224; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_226 = 8'he2 == inBytes_0 ? 8'h98 : _GEN_225; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_227 = 8'he3 == inBytes_0 ? 8'h11 : _GEN_226; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_228 = 8'he4 == inBytes_0 ? 8'h69 : _GEN_227; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_229 = 8'he5 == inBytes_0 ? 8'hd9 : _GEN_228; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_230 = 8'he6 == inBytes_0 ? 8'h8e : _GEN_229; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_231 = 8'he7 == inBytes_0 ? 8'h94 : _GEN_230; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_232 = 8'he8 == inBytes_0 ? 8'h9b : _GEN_231; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_233 = 8'he9 == inBytes_0 ? 8'h1e : _GEN_232; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_234 = 8'hea == inBytes_0 ? 8'h87 : _GEN_233; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_235 = 8'heb == inBytes_0 ? 8'he9 : _GEN_234; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_236 = 8'hec == inBytes_0 ? 8'hce : _GEN_235; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_237 = 8'hed == inBytes_0 ? 8'h55 : _GEN_236; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_238 = 8'hee == inBytes_0 ? 8'h28 : _GEN_237; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_239 = 8'hef == inBytes_0 ? 8'hdf : _GEN_238; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_240 = 8'hf0 == inBytes_0 ? 8'h8c : _GEN_239; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_241 = 8'hf1 == inBytes_0 ? 8'ha1 : _GEN_240; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_242 = 8'hf2 == inBytes_0 ? 8'h89 : _GEN_241; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_243 = 8'hf3 == inBytes_0 ? 8'hd : _GEN_242; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_244 = 8'hf4 == inBytes_0 ? 8'hbf : _GEN_243; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_245 = 8'hf5 == inBytes_0 ? 8'he6 : _GEN_244; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_246 = 8'hf6 == inBytes_0 ? 8'h42 : _GEN_245; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_247 = 8'hf7 == inBytes_0 ? 8'h68 : _GEN_246; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_248 = 8'hf8 == inBytes_0 ? 8'h41 : _GEN_247; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_249 = 8'hf9 == inBytes_0 ? 8'h99 : _GEN_248; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_250 = 8'hfa == inBytes_0 ? 8'h2d : _GEN_249; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_251 = 8'hfb == inBytes_0 ? 8'hf : _GEN_250; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_252 = 8'hfc == inBytes_0 ? 8'hb0 : _GEN_251; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_253 = 8'hfd == inBytes_0 ? 8'h54 : _GEN_252; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_254 = 8'hfe == inBytes_0 ? 8'hbb : _GEN_253; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] outBytes_0 = 8'hff == inBytes_0 ? 8'h16 : _GEN_254; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_257 = 8'h1 == inBytes_1 ? 8'h7c : 8'h63; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_258 = 8'h2 == inBytes_1 ? 8'h77 : _GEN_257; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_259 = 8'h3 == inBytes_1 ? 8'h7b : _GEN_258; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_260 = 8'h4 == inBytes_1 ? 8'hf2 : _GEN_259; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_261 = 8'h5 == inBytes_1 ? 8'h6b : _GEN_260; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_262 = 8'h6 == inBytes_1 ? 8'h6f : _GEN_261; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_263 = 8'h7 == inBytes_1 ? 8'hc5 : _GEN_262; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_264 = 8'h8 == inBytes_1 ? 8'h30 : _GEN_263; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_265 = 8'h9 == inBytes_1 ? 8'h1 : _GEN_264; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_266 = 8'ha == inBytes_1 ? 8'h67 : _GEN_265; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_267 = 8'hb == inBytes_1 ? 8'h2b : _GEN_266; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_268 = 8'hc == inBytes_1 ? 8'hfe : _GEN_267; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_269 = 8'hd == inBytes_1 ? 8'hd7 : _GEN_268; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_270 = 8'he == inBytes_1 ? 8'hab : _GEN_269; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_271 = 8'hf == inBytes_1 ? 8'h76 : _GEN_270; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_272 = 8'h10 == inBytes_1 ? 8'hca : _GEN_271; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_273 = 8'h11 == inBytes_1 ? 8'h82 : _GEN_272; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_274 = 8'h12 == inBytes_1 ? 8'hc9 : _GEN_273; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_275 = 8'h13 == inBytes_1 ? 8'h7d : _GEN_274; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_276 = 8'h14 == inBytes_1 ? 8'hfa : _GEN_275; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_277 = 8'h15 == inBytes_1 ? 8'h59 : _GEN_276; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_278 = 8'h16 == inBytes_1 ? 8'h47 : _GEN_277; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_279 = 8'h17 == inBytes_1 ? 8'hf0 : _GEN_278; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_280 = 8'h18 == inBytes_1 ? 8'had : _GEN_279; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_281 = 8'h19 == inBytes_1 ? 8'hd4 : _GEN_280; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_282 = 8'h1a == inBytes_1 ? 8'ha2 : _GEN_281; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_283 = 8'h1b == inBytes_1 ? 8'haf : _GEN_282; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_284 = 8'h1c == inBytes_1 ? 8'h9c : _GEN_283; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_285 = 8'h1d == inBytes_1 ? 8'ha4 : _GEN_284; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_286 = 8'h1e == inBytes_1 ? 8'h72 : _GEN_285; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_287 = 8'h1f == inBytes_1 ? 8'hc0 : _GEN_286; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_288 = 8'h20 == inBytes_1 ? 8'hb7 : _GEN_287; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_289 = 8'h21 == inBytes_1 ? 8'hfd : _GEN_288; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_290 = 8'h22 == inBytes_1 ? 8'h93 : _GEN_289; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_291 = 8'h23 == inBytes_1 ? 8'h26 : _GEN_290; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_292 = 8'h24 == inBytes_1 ? 8'h36 : _GEN_291; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_293 = 8'h25 == inBytes_1 ? 8'h3f : _GEN_292; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_294 = 8'h26 == inBytes_1 ? 8'hf7 : _GEN_293; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_295 = 8'h27 == inBytes_1 ? 8'hcc : _GEN_294; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_296 = 8'h28 == inBytes_1 ? 8'h34 : _GEN_295; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_297 = 8'h29 == inBytes_1 ? 8'ha5 : _GEN_296; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_298 = 8'h2a == inBytes_1 ? 8'he5 : _GEN_297; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_299 = 8'h2b == inBytes_1 ? 8'hf1 : _GEN_298; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_300 = 8'h2c == inBytes_1 ? 8'h71 : _GEN_299; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_301 = 8'h2d == inBytes_1 ? 8'hd8 : _GEN_300; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_302 = 8'h2e == inBytes_1 ? 8'h31 : _GEN_301; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_303 = 8'h2f == inBytes_1 ? 8'h15 : _GEN_302; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_304 = 8'h30 == inBytes_1 ? 8'h4 : _GEN_303; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_305 = 8'h31 == inBytes_1 ? 8'hc7 : _GEN_304; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_306 = 8'h32 == inBytes_1 ? 8'h23 : _GEN_305; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_307 = 8'h33 == inBytes_1 ? 8'hc3 : _GEN_306; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_308 = 8'h34 == inBytes_1 ? 8'h18 : _GEN_307; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_309 = 8'h35 == inBytes_1 ? 8'h96 : _GEN_308; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_310 = 8'h36 == inBytes_1 ? 8'h5 : _GEN_309; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_311 = 8'h37 == inBytes_1 ? 8'h9a : _GEN_310; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_312 = 8'h38 == inBytes_1 ? 8'h7 : _GEN_311; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_313 = 8'h39 == inBytes_1 ? 8'h12 : _GEN_312; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_314 = 8'h3a == inBytes_1 ? 8'h80 : _GEN_313; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_315 = 8'h3b == inBytes_1 ? 8'he2 : _GEN_314; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_316 = 8'h3c == inBytes_1 ? 8'heb : _GEN_315; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_317 = 8'h3d == inBytes_1 ? 8'h27 : _GEN_316; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_318 = 8'h3e == inBytes_1 ? 8'hb2 : _GEN_317; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_319 = 8'h3f == inBytes_1 ? 8'h75 : _GEN_318; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_320 = 8'h40 == inBytes_1 ? 8'h9 : _GEN_319; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_321 = 8'h41 == inBytes_1 ? 8'h83 : _GEN_320; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_322 = 8'h42 == inBytes_1 ? 8'h2c : _GEN_321; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_323 = 8'h43 == inBytes_1 ? 8'h1a : _GEN_322; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_324 = 8'h44 == inBytes_1 ? 8'h1b : _GEN_323; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_325 = 8'h45 == inBytes_1 ? 8'h6e : _GEN_324; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_326 = 8'h46 == inBytes_1 ? 8'h5a : _GEN_325; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_327 = 8'h47 == inBytes_1 ? 8'ha0 : _GEN_326; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_328 = 8'h48 == inBytes_1 ? 8'h52 : _GEN_327; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_329 = 8'h49 == inBytes_1 ? 8'h3b : _GEN_328; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_330 = 8'h4a == inBytes_1 ? 8'hd6 : _GEN_329; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_331 = 8'h4b == inBytes_1 ? 8'hb3 : _GEN_330; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_332 = 8'h4c == inBytes_1 ? 8'h29 : _GEN_331; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_333 = 8'h4d == inBytes_1 ? 8'he3 : _GEN_332; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_334 = 8'h4e == inBytes_1 ? 8'h2f : _GEN_333; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_335 = 8'h4f == inBytes_1 ? 8'h84 : _GEN_334; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_336 = 8'h50 == inBytes_1 ? 8'h53 : _GEN_335; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_337 = 8'h51 == inBytes_1 ? 8'hd1 : _GEN_336; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_338 = 8'h52 == inBytes_1 ? 8'h0 : _GEN_337; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_339 = 8'h53 == inBytes_1 ? 8'hed : _GEN_338; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_340 = 8'h54 == inBytes_1 ? 8'h20 : _GEN_339; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_341 = 8'h55 == inBytes_1 ? 8'hfc : _GEN_340; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_342 = 8'h56 == inBytes_1 ? 8'hb1 : _GEN_341; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_343 = 8'h57 == inBytes_1 ? 8'h5b : _GEN_342; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_344 = 8'h58 == inBytes_1 ? 8'h6a : _GEN_343; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_345 = 8'h59 == inBytes_1 ? 8'hcb : _GEN_344; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_346 = 8'h5a == inBytes_1 ? 8'hbe : _GEN_345; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_347 = 8'h5b == inBytes_1 ? 8'h39 : _GEN_346; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_348 = 8'h5c == inBytes_1 ? 8'h4a : _GEN_347; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_349 = 8'h5d == inBytes_1 ? 8'h4c : _GEN_348; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_350 = 8'h5e == inBytes_1 ? 8'h58 : _GEN_349; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_351 = 8'h5f == inBytes_1 ? 8'hcf : _GEN_350; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_352 = 8'h60 == inBytes_1 ? 8'hd0 : _GEN_351; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_353 = 8'h61 == inBytes_1 ? 8'hef : _GEN_352; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_354 = 8'h62 == inBytes_1 ? 8'haa : _GEN_353; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_355 = 8'h63 == inBytes_1 ? 8'hfb : _GEN_354; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_356 = 8'h64 == inBytes_1 ? 8'h43 : _GEN_355; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_357 = 8'h65 == inBytes_1 ? 8'h4d : _GEN_356; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_358 = 8'h66 == inBytes_1 ? 8'h33 : _GEN_357; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_359 = 8'h67 == inBytes_1 ? 8'h85 : _GEN_358; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_360 = 8'h68 == inBytes_1 ? 8'h45 : _GEN_359; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_361 = 8'h69 == inBytes_1 ? 8'hf9 : _GEN_360; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_362 = 8'h6a == inBytes_1 ? 8'h2 : _GEN_361; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_363 = 8'h6b == inBytes_1 ? 8'h7f : _GEN_362; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_364 = 8'h6c == inBytes_1 ? 8'h50 : _GEN_363; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_365 = 8'h6d == inBytes_1 ? 8'h3c : _GEN_364; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_366 = 8'h6e == inBytes_1 ? 8'h9f : _GEN_365; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_367 = 8'h6f == inBytes_1 ? 8'ha8 : _GEN_366; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_368 = 8'h70 == inBytes_1 ? 8'h51 : _GEN_367; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_369 = 8'h71 == inBytes_1 ? 8'ha3 : _GEN_368; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_370 = 8'h72 == inBytes_1 ? 8'h40 : _GEN_369; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_371 = 8'h73 == inBytes_1 ? 8'h8f : _GEN_370; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_372 = 8'h74 == inBytes_1 ? 8'h92 : _GEN_371; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_373 = 8'h75 == inBytes_1 ? 8'h9d : _GEN_372; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_374 = 8'h76 == inBytes_1 ? 8'h38 : _GEN_373; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_375 = 8'h77 == inBytes_1 ? 8'hf5 : _GEN_374; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_376 = 8'h78 == inBytes_1 ? 8'hbc : _GEN_375; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_377 = 8'h79 == inBytes_1 ? 8'hb6 : _GEN_376; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_378 = 8'h7a == inBytes_1 ? 8'hda : _GEN_377; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_379 = 8'h7b == inBytes_1 ? 8'h21 : _GEN_378; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_380 = 8'h7c == inBytes_1 ? 8'h10 : _GEN_379; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_381 = 8'h7d == inBytes_1 ? 8'hff : _GEN_380; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_382 = 8'h7e == inBytes_1 ? 8'hf3 : _GEN_381; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_383 = 8'h7f == inBytes_1 ? 8'hd2 : _GEN_382; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_384 = 8'h80 == inBytes_1 ? 8'hcd : _GEN_383; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_385 = 8'h81 == inBytes_1 ? 8'hc : _GEN_384; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_386 = 8'h82 == inBytes_1 ? 8'h13 : _GEN_385; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_387 = 8'h83 == inBytes_1 ? 8'hec : _GEN_386; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_388 = 8'h84 == inBytes_1 ? 8'h5f : _GEN_387; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_389 = 8'h85 == inBytes_1 ? 8'h97 : _GEN_388; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_390 = 8'h86 == inBytes_1 ? 8'h44 : _GEN_389; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_391 = 8'h87 == inBytes_1 ? 8'h17 : _GEN_390; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_392 = 8'h88 == inBytes_1 ? 8'hc4 : _GEN_391; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_393 = 8'h89 == inBytes_1 ? 8'ha7 : _GEN_392; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_394 = 8'h8a == inBytes_1 ? 8'h7e : _GEN_393; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_395 = 8'h8b == inBytes_1 ? 8'h3d : _GEN_394; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_396 = 8'h8c == inBytes_1 ? 8'h64 : _GEN_395; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_397 = 8'h8d == inBytes_1 ? 8'h5d : _GEN_396; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_398 = 8'h8e == inBytes_1 ? 8'h19 : _GEN_397; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_399 = 8'h8f == inBytes_1 ? 8'h73 : _GEN_398; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_400 = 8'h90 == inBytes_1 ? 8'h60 : _GEN_399; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_401 = 8'h91 == inBytes_1 ? 8'h81 : _GEN_400; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_402 = 8'h92 == inBytes_1 ? 8'h4f : _GEN_401; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_403 = 8'h93 == inBytes_1 ? 8'hdc : _GEN_402; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_404 = 8'h94 == inBytes_1 ? 8'h22 : _GEN_403; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_405 = 8'h95 == inBytes_1 ? 8'h2a : _GEN_404; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_406 = 8'h96 == inBytes_1 ? 8'h90 : _GEN_405; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_407 = 8'h97 == inBytes_1 ? 8'h88 : _GEN_406; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_408 = 8'h98 == inBytes_1 ? 8'h46 : _GEN_407; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_409 = 8'h99 == inBytes_1 ? 8'hee : _GEN_408; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_410 = 8'h9a == inBytes_1 ? 8'hb8 : _GEN_409; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_411 = 8'h9b == inBytes_1 ? 8'h14 : _GEN_410; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_412 = 8'h9c == inBytes_1 ? 8'hde : _GEN_411; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_413 = 8'h9d == inBytes_1 ? 8'h5e : _GEN_412; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_414 = 8'h9e == inBytes_1 ? 8'hb : _GEN_413; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_415 = 8'h9f == inBytes_1 ? 8'hdb : _GEN_414; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_416 = 8'ha0 == inBytes_1 ? 8'he0 : _GEN_415; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_417 = 8'ha1 == inBytes_1 ? 8'h32 : _GEN_416; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_418 = 8'ha2 == inBytes_1 ? 8'h3a : _GEN_417; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_419 = 8'ha3 == inBytes_1 ? 8'ha : _GEN_418; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_420 = 8'ha4 == inBytes_1 ? 8'h49 : _GEN_419; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_421 = 8'ha5 == inBytes_1 ? 8'h6 : _GEN_420; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_422 = 8'ha6 == inBytes_1 ? 8'h24 : _GEN_421; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_423 = 8'ha7 == inBytes_1 ? 8'h5c : _GEN_422; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_424 = 8'ha8 == inBytes_1 ? 8'hc2 : _GEN_423; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_425 = 8'ha9 == inBytes_1 ? 8'hd3 : _GEN_424; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_426 = 8'haa == inBytes_1 ? 8'hac : _GEN_425; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_427 = 8'hab == inBytes_1 ? 8'h62 : _GEN_426; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_428 = 8'hac == inBytes_1 ? 8'h91 : _GEN_427; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_429 = 8'had == inBytes_1 ? 8'h95 : _GEN_428; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_430 = 8'hae == inBytes_1 ? 8'he4 : _GEN_429; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_431 = 8'haf == inBytes_1 ? 8'h79 : _GEN_430; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_432 = 8'hb0 == inBytes_1 ? 8'he7 : _GEN_431; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_433 = 8'hb1 == inBytes_1 ? 8'hc8 : _GEN_432; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_434 = 8'hb2 == inBytes_1 ? 8'h37 : _GEN_433; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_435 = 8'hb3 == inBytes_1 ? 8'h6d : _GEN_434; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_436 = 8'hb4 == inBytes_1 ? 8'h8d : _GEN_435; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_437 = 8'hb5 == inBytes_1 ? 8'hd5 : _GEN_436; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_438 = 8'hb6 == inBytes_1 ? 8'h4e : _GEN_437; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_439 = 8'hb7 == inBytes_1 ? 8'ha9 : _GEN_438; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_440 = 8'hb8 == inBytes_1 ? 8'h6c : _GEN_439; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_441 = 8'hb9 == inBytes_1 ? 8'h56 : _GEN_440; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_442 = 8'hba == inBytes_1 ? 8'hf4 : _GEN_441; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_443 = 8'hbb == inBytes_1 ? 8'hea : _GEN_442; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_444 = 8'hbc == inBytes_1 ? 8'h65 : _GEN_443; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_445 = 8'hbd == inBytes_1 ? 8'h7a : _GEN_444; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_446 = 8'hbe == inBytes_1 ? 8'hae : _GEN_445; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_447 = 8'hbf == inBytes_1 ? 8'h8 : _GEN_446; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_448 = 8'hc0 == inBytes_1 ? 8'hba : _GEN_447; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_449 = 8'hc1 == inBytes_1 ? 8'h78 : _GEN_448; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_450 = 8'hc2 == inBytes_1 ? 8'h25 : _GEN_449; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_451 = 8'hc3 == inBytes_1 ? 8'h2e : _GEN_450; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_452 = 8'hc4 == inBytes_1 ? 8'h1c : _GEN_451; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_453 = 8'hc5 == inBytes_1 ? 8'ha6 : _GEN_452; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_454 = 8'hc6 == inBytes_1 ? 8'hb4 : _GEN_453; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_455 = 8'hc7 == inBytes_1 ? 8'hc6 : _GEN_454; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_456 = 8'hc8 == inBytes_1 ? 8'he8 : _GEN_455; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_457 = 8'hc9 == inBytes_1 ? 8'hdd : _GEN_456; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_458 = 8'hca == inBytes_1 ? 8'h74 : _GEN_457; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_459 = 8'hcb == inBytes_1 ? 8'h1f : _GEN_458; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_460 = 8'hcc == inBytes_1 ? 8'h4b : _GEN_459; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_461 = 8'hcd == inBytes_1 ? 8'hbd : _GEN_460; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_462 = 8'hce == inBytes_1 ? 8'h8b : _GEN_461; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_463 = 8'hcf == inBytes_1 ? 8'h8a : _GEN_462; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_464 = 8'hd0 == inBytes_1 ? 8'h70 : _GEN_463; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_465 = 8'hd1 == inBytes_1 ? 8'h3e : _GEN_464; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_466 = 8'hd2 == inBytes_1 ? 8'hb5 : _GEN_465; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_467 = 8'hd3 == inBytes_1 ? 8'h66 : _GEN_466; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_468 = 8'hd4 == inBytes_1 ? 8'h48 : _GEN_467; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_469 = 8'hd5 == inBytes_1 ? 8'h3 : _GEN_468; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_470 = 8'hd6 == inBytes_1 ? 8'hf6 : _GEN_469; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_471 = 8'hd7 == inBytes_1 ? 8'he : _GEN_470; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_472 = 8'hd8 == inBytes_1 ? 8'h61 : _GEN_471; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_473 = 8'hd9 == inBytes_1 ? 8'h35 : _GEN_472; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_474 = 8'hda == inBytes_1 ? 8'h57 : _GEN_473; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_475 = 8'hdb == inBytes_1 ? 8'hb9 : _GEN_474; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_476 = 8'hdc == inBytes_1 ? 8'h86 : _GEN_475; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_477 = 8'hdd == inBytes_1 ? 8'hc1 : _GEN_476; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_478 = 8'hde == inBytes_1 ? 8'h1d : _GEN_477; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_479 = 8'hdf == inBytes_1 ? 8'h9e : _GEN_478; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_480 = 8'he0 == inBytes_1 ? 8'he1 : _GEN_479; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_481 = 8'he1 == inBytes_1 ? 8'hf8 : _GEN_480; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_482 = 8'he2 == inBytes_1 ? 8'h98 : _GEN_481; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_483 = 8'he3 == inBytes_1 ? 8'h11 : _GEN_482; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_484 = 8'he4 == inBytes_1 ? 8'h69 : _GEN_483; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_485 = 8'he5 == inBytes_1 ? 8'hd9 : _GEN_484; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_486 = 8'he6 == inBytes_1 ? 8'h8e : _GEN_485; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_487 = 8'he7 == inBytes_1 ? 8'h94 : _GEN_486; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_488 = 8'he8 == inBytes_1 ? 8'h9b : _GEN_487; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_489 = 8'he9 == inBytes_1 ? 8'h1e : _GEN_488; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_490 = 8'hea == inBytes_1 ? 8'h87 : _GEN_489; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_491 = 8'heb == inBytes_1 ? 8'he9 : _GEN_490; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_492 = 8'hec == inBytes_1 ? 8'hce : _GEN_491; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_493 = 8'hed == inBytes_1 ? 8'h55 : _GEN_492; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_494 = 8'hee == inBytes_1 ? 8'h28 : _GEN_493; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_495 = 8'hef == inBytes_1 ? 8'hdf : _GEN_494; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_496 = 8'hf0 == inBytes_1 ? 8'h8c : _GEN_495; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_497 = 8'hf1 == inBytes_1 ? 8'ha1 : _GEN_496; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_498 = 8'hf2 == inBytes_1 ? 8'h89 : _GEN_497; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_499 = 8'hf3 == inBytes_1 ? 8'hd : _GEN_498; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_500 = 8'hf4 == inBytes_1 ? 8'hbf : _GEN_499; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_501 = 8'hf5 == inBytes_1 ? 8'he6 : _GEN_500; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_502 = 8'hf6 == inBytes_1 ? 8'h42 : _GEN_501; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_503 = 8'hf7 == inBytes_1 ? 8'h68 : _GEN_502; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_504 = 8'hf8 == inBytes_1 ? 8'h41 : _GEN_503; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_505 = 8'hf9 == inBytes_1 ? 8'h99 : _GEN_504; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_506 = 8'hfa == inBytes_1 ? 8'h2d : _GEN_505; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_507 = 8'hfb == inBytes_1 ? 8'hf : _GEN_506; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_508 = 8'hfc == inBytes_1 ? 8'hb0 : _GEN_507; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_509 = 8'hfd == inBytes_1 ? 8'h54 : _GEN_508; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_510 = 8'hfe == inBytes_1 ? 8'hbb : _GEN_509; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] outBytes_1 = 8'hff == inBytes_1 ? 8'h16 : _GEN_510; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_513 = 8'h1 == inBytes_2 ? 8'h7c : 8'h63; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_514 = 8'h2 == inBytes_2 ? 8'h77 : _GEN_513; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_515 = 8'h3 == inBytes_2 ? 8'h7b : _GEN_514; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_516 = 8'h4 == inBytes_2 ? 8'hf2 : _GEN_515; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_517 = 8'h5 == inBytes_2 ? 8'h6b : _GEN_516; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_518 = 8'h6 == inBytes_2 ? 8'h6f : _GEN_517; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_519 = 8'h7 == inBytes_2 ? 8'hc5 : _GEN_518; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_520 = 8'h8 == inBytes_2 ? 8'h30 : _GEN_519; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_521 = 8'h9 == inBytes_2 ? 8'h1 : _GEN_520; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_522 = 8'ha == inBytes_2 ? 8'h67 : _GEN_521; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_523 = 8'hb == inBytes_2 ? 8'h2b : _GEN_522; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_524 = 8'hc == inBytes_2 ? 8'hfe : _GEN_523; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_525 = 8'hd == inBytes_2 ? 8'hd7 : _GEN_524; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_526 = 8'he == inBytes_2 ? 8'hab : _GEN_525; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_527 = 8'hf == inBytes_2 ? 8'h76 : _GEN_526; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_528 = 8'h10 == inBytes_2 ? 8'hca : _GEN_527; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_529 = 8'h11 == inBytes_2 ? 8'h82 : _GEN_528; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_530 = 8'h12 == inBytes_2 ? 8'hc9 : _GEN_529; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_531 = 8'h13 == inBytes_2 ? 8'h7d : _GEN_530; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_532 = 8'h14 == inBytes_2 ? 8'hfa : _GEN_531; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_533 = 8'h15 == inBytes_2 ? 8'h59 : _GEN_532; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_534 = 8'h16 == inBytes_2 ? 8'h47 : _GEN_533; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_535 = 8'h17 == inBytes_2 ? 8'hf0 : _GEN_534; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_536 = 8'h18 == inBytes_2 ? 8'had : _GEN_535; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_537 = 8'h19 == inBytes_2 ? 8'hd4 : _GEN_536; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_538 = 8'h1a == inBytes_2 ? 8'ha2 : _GEN_537; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_539 = 8'h1b == inBytes_2 ? 8'haf : _GEN_538; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_540 = 8'h1c == inBytes_2 ? 8'h9c : _GEN_539; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_541 = 8'h1d == inBytes_2 ? 8'ha4 : _GEN_540; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_542 = 8'h1e == inBytes_2 ? 8'h72 : _GEN_541; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_543 = 8'h1f == inBytes_2 ? 8'hc0 : _GEN_542; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_544 = 8'h20 == inBytes_2 ? 8'hb7 : _GEN_543; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_545 = 8'h21 == inBytes_2 ? 8'hfd : _GEN_544; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_546 = 8'h22 == inBytes_2 ? 8'h93 : _GEN_545; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_547 = 8'h23 == inBytes_2 ? 8'h26 : _GEN_546; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_548 = 8'h24 == inBytes_2 ? 8'h36 : _GEN_547; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_549 = 8'h25 == inBytes_2 ? 8'h3f : _GEN_548; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_550 = 8'h26 == inBytes_2 ? 8'hf7 : _GEN_549; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_551 = 8'h27 == inBytes_2 ? 8'hcc : _GEN_550; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_552 = 8'h28 == inBytes_2 ? 8'h34 : _GEN_551; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_553 = 8'h29 == inBytes_2 ? 8'ha5 : _GEN_552; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_554 = 8'h2a == inBytes_2 ? 8'he5 : _GEN_553; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_555 = 8'h2b == inBytes_2 ? 8'hf1 : _GEN_554; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_556 = 8'h2c == inBytes_2 ? 8'h71 : _GEN_555; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_557 = 8'h2d == inBytes_2 ? 8'hd8 : _GEN_556; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_558 = 8'h2e == inBytes_2 ? 8'h31 : _GEN_557; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_559 = 8'h2f == inBytes_2 ? 8'h15 : _GEN_558; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_560 = 8'h30 == inBytes_2 ? 8'h4 : _GEN_559; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_561 = 8'h31 == inBytes_2 ? 8'hc7 : _GEN_560; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_562 = 8'h32 == inBytes_2 ? 8'h23 : _GEN_561; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_563 = 8'h33 == inBytes_2 ? 8'hc3 : _GEN_562; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_564 = 8'h34 == inBytes_2 ? 8'h18 : _GEN_563; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_565 = 8'h35 == inBytes_2 ? 8'h96 : _GEN_564; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_566 = 8'h36 == inBytes_2 ? 8'h5 : _GEN_565; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_567 = 8'h37 == inBytes_2 ? 8'h9a : _GEN_566; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_568 = 8'h38 == inBytes_2 ? 8'h7 : _GEN_567; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_569 = 8'h39 == inBytes_2 ? 8'h12 : _GEN_568; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_570 = 8'h3a == inBytes_2 ? 8'h80 : _GEN_569; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_571 = 8'h3b == inBytes_2 ? 8'he2 : _GEN_570; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_572 = 8'h3c == inBytes_2 ? 8'heb : _GEN_571; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_573 = 8'h3d == inBytes_2 ? 8'h27 : _GEN_572; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_574 = 8'h3e == inBytes_2 ? 8'hb2 : _GEN_573; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_575 = 8'h3f == inBytes_2 ? 8'h75 : _GEN_574; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_576 = 8'h40 == inBytes_2 ? 8'h9 : _GEN_575; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_577 = 8'h41 == inBytes_2 ? 8'h83 : _GEN_576; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_578 = 8'h42 == inBytes_2 ? 8'h2c : _GEN_577; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_579 = 8'h43 == inBytes_2 ? 8'h1a : _GEN_578; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_580 = 8'h44 == inBytes_2 ? 8'h1b : _GEN_579; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_581 = 8'h45 == inBytes_2 ? 8'h6e : _GEN_580; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_582 = 8'h46 == inBytes_2 ? 8'h5a : _GEN_581; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_583 = 8'h47 == inBytes_2 ? 8'ha0 : _GEN_582; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_584 = 8'h48 == inBytes_2 ? 8'h52 : _GEN_583; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_585 = 8'h49 == inBytes_2 ? 8'h3b : _GEN_584; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_586 = 8'h4a == inBytes_2 ? 8'hd6 : _GEN_585; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_587 = 8'h4b == inBytes_2 ? 8'hb3 : _GEN_586; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_588 = 8'h4c == inBytes_2 ? 8'h29 : _GEN_587; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_589 = 8'h4d == inBytes_2 ? 8'he3 : _GEN_588; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_590 = 8'h4e == inBytes_2 ? 8'h2f : _GEN_589; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_591 = 8'h4f == inBytes_2 ? 8'h84 : _GEN_590; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_592 = 8'h50 == inBytes_2 ? 8'h53 : _GEN_591; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_593 = 8'h51 == inBytes_2 ? 8'hd1 : _GEN_592; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_594 = 8'h52 == inBytes_2 ? 8'h0 : _GEN_593; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_595 = 8'h53 == inBytes_2 ? 8'hed : _GEN_594; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_596 = 8'h54 == inBytes_2 ? 8'h20 : _GEN_595; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_597 = 8'h55 == inBytes_2 ? 8'hfc : _GEN_596; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_598 = 8'h56 == inBytes_2 ? 8'hb1 : _GEN_597; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_599 = 8'h57 == inBytes_2 ? 8'h5b : _GEN_598; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_600 = 8'h58 == inBytes_2 ? 8'h6a : _GEN_599; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_601 = 8'h59 == inBytes_2 ? 8'hcb : _GEN_600; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_602 = 8'h5a == inBytes_2 ? 8'hbe : _GEN_601; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_603 = 8'h5b == inBytes_2 ? 8'h39 : _GEN_602; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_604 = 8'h5c == inBytes_2 ? 8'h4a : _GEN_603; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_605 = 8'h5d == inBytes_2 ? 8'h4c : _GEN_604; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_606 = 8'h5e == inBytes_2 ? 8'h58 : _GEN_605; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_607 = 8'h5f == inBytes_2 ? 8'hcf : _GEN_606; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_608 = 8'h60 == inBytes_2 ? 8'hd0 : _GEN_607; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_609 = 8'h61 == inBytes_2 ? 8'hef : _GEN_608; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_610 = 8'h62 == inBytes_2 ? 8'haa : _GEN_609; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_611 = 8'h63 == inBytes_2 ? 8'hfb : _GEN_610; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_612 = 8'h64 == inBytes_2 ? 8'h43 : _GEN_611; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_613 = 8'h65 == inBytes_2 ? 8'h4d : _GEN_612; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_614 = 8'h66 == inBytes_2 ? 8'h33 : _GEN_613; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_615 = 8'h67 == inBytes_2 ? 8'h85 : _GEN_614; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_616 = 8'h68 == inBytes_2 ? 8'h45 : _GEN_615; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_617 = 8'h69 == inBytes_2 ? 8'hf9 : _GEN_616; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_618 = 8'h6a == inBytes_2 ? 8'h2 : _GEN_617; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_619 = 8'h6b == inBytes_2 ? 8'h7f : _GEN_618; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_620 = 8'h6c == inBytes_2 ? 8'h50 : _GEN_619; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_621 = 8'h6d == inBytes_2 ? 8'h3c : _GEN_620; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_622 = 8'h6e == inBytes_2 ? 8'h9f : _GEN_621; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_623 = 8'h6f == inBytes_2 ? 8'ha8 : _GEN_622; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_624 = 8'h70 == inBytes_2 ? 8'h51 : _GEN_623; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_625 = 8'h71 == inBytes_2 ? 8'ha3 : _GEN_624; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_626 = 8'h72 == inBytes_2 ? 8'h40 : _GEN_625; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_627 = 8'h73 == inBytes_2 ? 8'h8f : _GEN_626; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_628 = 8'h74 == inBytes_2 ? 8'h92 : _GEN_627; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_629 = 8'h75 == inBytes_2 ? 8'h9d : _GEN_628; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_630 = 8'h76 == inBytes_2 ? 8'h38 : _GEN_629; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_631 = 8'h77 == inBytes_2 ? 8'hf5 : _GEN_630; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_632 = 8'h78 == inBytes_2 ? 8'hbc : _GEN_631; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_633 = 8'h79 == inBytes_2 ? 8'hb6 : _GEN_632; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_634 = 8'h7a == inBytes_2 ? 8'hda : _GEN_633; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_635 = 8'h7b == inBytes_2 ? 8'h21 : _GEN_634; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_636 = 8'h7c == inBytes_2 ? 8'h10 : _GEN_635; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_637 = 8'h7d == inBytes_2 ? 8'hff : _GEN_636; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_638 = 8'h7e == inBytes_2 ? 8'hf3 : _GEN_637; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_639 = 8'h7f == inBytes_2 ? 8'hd2 : _GEN_638; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_640 = 8'h80 == inBytes_2 ? 8'hcd : _GEN_639; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_641 = 8'h81 == inBytes_2 ? 8'hc : _GEN_640; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_642 = 8'h82 == inBytes_2 ? 8'h13 : _GEN_641; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_643 = 8'h83 == inBytes_2 ? 8'hec : _GEN_642; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_644 = 8'h84 == inBytes_2 ? 8'h5f : _GEN_643; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_645 = 8'h85 == inBytes_2 ? 8'h97 : _GEN_644; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_646 = 8'h86 == inBytes_2 ? 8'h44 : _GEN_645; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_647 = 8'h87 == inBytes_2 ? 8'h17 : _GEN_646; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_648 = 8'h88 == inBytes_2 ? 8'hc4 : _GEN_647; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_649 = 8'h89 == inBytes_2 ? 8'ha7 : _GEN_648; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_650 = 8'h8a == inBytes_2 ? 8'h7e : _GEN_649; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_651 = 8'h8b == inBytes_2 ? 8'h3d : _GEN_650; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_652 = 8'h8c == inBytes_2 ? 8'h64 : _GEN_651; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_653 = 8'h8d == inBytes_2 ? 8'h5d : _GEN_652; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_654 = 8'h8e == inBytes_2 ? 8'h19 : _GEN_653; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_655 = 8'h8f == inBytes_2 ? 8'h73 : _GEN_654; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_656 = 8'h90 == inBytes_2 ? 8'h60 : _GEN_655; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_657 = 8'h91 == inBytes_2 ? 8'h81 : _GEN_656; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_658 = 8'h92 == inBytes_2 ? 8'h4f : _GEN_657; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_659 = 8'h93 == inBytes_2 ? 8'hdc : _GEN_658; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_660 = 8'h94 == inBytes_2 ? 8'h22 : _GEN_659; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_661 = 8'h95 == inBytes_2 ? 8'h2a : _GEN_660; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_662 = 8'h96 == inBytes_2 ? 8'h90 : _GEN_661; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_663 = 8'h97 == inBytes_2 ? 8'h88 : _GEN_662; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_664 = 8'h98 == inBytes_2 ? 8'h46 : _GEN_663; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_665 = 8'h99 == inBytes_2 ? 8'hee : _GEN_664; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_666 = 8'h9a == inBytes_2 ? 8'hb8 : _GEN_665; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_667 = 8'h9b == inBytes_2 ? 8'h14 : _GEN_666; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_668 = 8'h9c == inBytes_2 ? 8'hde : _GEN_667; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_669 = 8'h9d == inBytes_2 ? 8'h5e : _GEN_668; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_670 = 8'h9e == inBytes_2 ? 8'hb : _GEN_669; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_671 = 8'h9f == inBytes_2 ? 8'hdb : _GEN_670; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_672 = 8'ha0 == inBytes_2 ? 8'he0 : _GEN_671; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_673 = 8'ha1 == inBytes_2 ? 8'h32 : _GEN_672; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_674 = 8'ha2 == inBytes_2 ? 8'h3a : _GEN_673; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_675 = 8'ha3 == inBytes_2 ? 8'ha : _GEN_674; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_676 = 8'ha4 == inBytes_2 ? 8'h49 : _GEN_675; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_677 = 8'ha5 == inBytes_2 ? 8'h6 : _GEN_676; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_678 = 8'ha6 == inBytes_2 ? 8'h24 : _GEN_677; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_679 = 8'ha7 == inBytes_2 ? 8'h5c : _GEN_678; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_680 = 8'ha8 == inBytes_2 ? 8'hc2 : _GEN_679; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_681 = 8'ha9 == inBytes_2 ? 8'hd3 : _GEN_680; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_682 = 8'haa == inBytes_2 ? 8'hac : _GEN_681; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_683 = 8'hab == inBytes_2 ? 8'h62 : _GEN_682; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_684 = 8'hac == inBytes_2 ? 8'h91 : _GEN_683; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_685 = 8'had == inBytes_2 ? 8'h95 : _GEN_684; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_686 = 8'hae == inBytes_2 ? 8'he4 : _GEN_685; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_687 = 8'haf == inBytes_2 ? 8'h79 : _GEN_686; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_688 = 8'hb0 == inBytes_2 ? 8'he7 : _GEN_687; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_689 = 8'hb1 == inBytes_2 ? 8'hc8 : _GEN_688; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_690 = 8'hb2 == inBytes_2 ? 8'h37 : _GEN_689; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_691 = 8'hb3 == inBytes_2 ? 8'h6d : _GEN_690; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_692 = 8'hb4 == inBytes_2 ? 8'h8d : _GEN_691; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_693 = 8'hb5 == inBytes_2 ? 8'hd5 : _GEN_692; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_694 = 8'hb6 == inBytes_2 ? 8'h4e : _GEN_693; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_695 = 8'hb7 == inBytes_2 ? 8'ha9 : _GEN_694; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_696 = 8'hb8 == inBytes_2 ? 8'h6c : _GEN_695; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_697 = 8'hb9 == inBytes_2 ? 8'h56 : _GEN_696; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_698 = 8'hba == inBytes_2 ? 8'hf4 : _GEN_697; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_699 = 8'hbb == inBytes_2 ? 8'hea : _GEN_698; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_700 = 8'hbc == inBytes_2 ? 8'h65 : _GEN_699; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_701 = 8'hbd == inBytes_2 ? 8'h7a : _GEN_700; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_702 = 8'hbe == inBytes_2 ? 8'hae : _GEN_701; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_703 = 8'hbf == inBytes_2 ? 8'h8 : _GEN_702; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_704 = 8'hc0 == inBytes_2 ? 8'hba : _GEN_703; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_705 = 8'hc1 == inBytes_2 ? 8'h78 : _GEN_704; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_706 = 8'hc2 == inBytes_2 ? 8'h25 : _GEN_705; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_707 = 8'hc3 == inBytes_2 ? 8'h2e : _GEN_706; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_708 = 8'hc4 == inBytes_2 ? 8'h1c : _GEN_707; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_709 = 8'hc5 == inBytes_2 ? 8'ha6 : _GEN_708; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_710 = 8'hc6 == inBytes_2 ? 8'hb4 : _GEN_709; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_711 = 8'hc7 == inBytes_2 ? 8'hc6 : _GEN_710; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_712 = 8'hc8 == inBytes_2 ? 8'he8 : _GEN_711; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_713 = 8'hc9 == inBytes_2 ? 8'hdd : _GEN_712; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_714 = 8'hca == inBytes_2 ? 8'h74 : _GEN_713; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_715 = 8'hcb == inBytes_2 ? 8'h1f : _GEN_714; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_716 = 8'hcc == inBytes_2 ? 8'h4b : _GEN_715; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_717 = 8'hcd == inBytes_2 ? 8'hbd : _GEN_716; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_718 = 8'hce == inBytes_2 ? 8'h8b : _GEN_717; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_719 = 8'hcf == inBytes_2 ? 8'h8a : _GEN_718; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_720 = 8'hd0 == inBytes_2 ? 8'h70 : _GEN_719; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_721 = 8'hd1 == inBytes_2 ? 8'h3e : _GEN_720; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_722 = 8'hd2 == inBytes_2 ? 8'hb5 : _GEN_721; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_723 = 8'hd3 == inBytes_2 ? 8'h66 : _GEN_722; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_724 = 8'hd4 == inBytes_2 ? 8'h48 : _GEN_723; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_725 = 8'hd5 == inBytes_2 ? 8'h3 : _GEN_724; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_726 = 8'hd6 == inBytes_2 ? 8'hf6 : _GEN_725; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_727 = 8'hd7 == inBytes_2 ? 8'he : _GEN_726; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_728 = 8'hd8 == inBytes_2 ? 8'h61 : _GEN_727; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_729 = 8'hd9 == inBytes_2 ? 8'h35 : _GEN_728; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_730 = 8'hda == inBytes_2 ? 8'h57 : _GEN_729; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_731 = 8'hdb == inBytes_2 ? 8'hb9 : _GEN_730; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_732 = 8'hdc == inBytes_2 ? 8'h86 : _GEN_731; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_733 = 8'hdd == inBytes_2 ? 8'hc1 : _GEN_732; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_734 = 8'hde == inBytes_2 ? 8'h1d : _GEN_733; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_735 = 8'hdf == inBytes_2 ? 8'h9e : _GEN_734; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_736 = 8'he0 == inBytes_2 ? 8'he1 : _GEN_735; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_737 = 8'he1 == inBytes_2 ? 8'hf8 : _GEN_736; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_738 = 8'he2 == inBytes_2 ? 8'h98 : _GEN_737; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_739 = 8'he3 == inBytes_2 ? 8'h11 : _GEN_738; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_740 = 8'he4 == inBytes_2 ? 8'h69 : _GEN_739; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_741 = 8'he5 == inBytes_2 ? 8'hd9 : _GEN_740; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_742 = 8'he6 == inBytes_2 ? 8'h8e : _GEN_741; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_743 = 8'he7 == inBytes_2 ? 8'h94 : _GEN_742; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_744 = 8'he8 == inBytes_2 ? 8'h9b : _GEN_743; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_745 = 8'he9 == inBytes_2 ? 8'h1e : _GEN_744; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_746 = 8'hea == inBytes_2 ? 8'h87 : _GEN_745; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_747 = 8'heb == inBytes_2 ? 8'he9 : _GEN_746; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_748 = 8'hec == inBytes_2 ? 8'hce : _GEN_747; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_749 = 8'hed == inBytes_2 ? 8'h55 : _GEN_748; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_750 = 8'hee == inBytes_2 ? 8'h28 : _GEN_749; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_751 = 8'hef == inBytes_2 ? 8'hdf : _GEN_750; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_752 = 8'hf0 == inBytes_2 ? 8'h8c : _GEN_751; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_753 = 8'hf1 == inBytes_2 ? 8'ha1 : _GEN_752; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_754 = 8'hf2 == inBytes_2 ? 8'h89 : _GEN_753; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_755 = 8'hf3 == inBytes_2 ? 8'hd : _GEN_754; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_756 = 8'hf4 == inBytes_2 ? 8'hbf : _GEN_755; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_757 = 8'hf5 == inBytes_2 ? 8'he6 : _GEN_756; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_758 = 8'hf6 == inBytes_2 ? 8'h42 : _GEN_757; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_759 = 8'hf7 == inBytes_2 ? 8'h68 : _GEN_758; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_760 = 8'hf8 == inBytes_2 ? 8'h41 : _GEN_759; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_761 = 8'hf9 == inBytes_2 ? 8'h99 : _GEN_760; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_762 = 8'hfa == inBytes_2 ? 8'h2d : _GEN_761; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_763 = 8'hfb == inBytes_2 ? 8'hf : _GEN_762; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_764 = 8'hfc == inBytes_2 ? 8'hb0 : _GEN_763; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_765 = 8'hfd == inBytes_2 ? 8'h54 : _GEN_764; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_766 = 8'hfe == inBytes_2 ? 8'hbb : _GEN_765; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] outBytes_2 = 8'hff == inBytes_2 ? 8'h16 : _GEN_766; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_769 = 8'h1 == inBytes_3 ? 8'h7c : 8'h63; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_770 = 8'h2 == inBytes_3 ? 8'h77 : _GEN_769; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_771 = 8'h3 == inBytes_3 ? 8'h7b : _GEN_770; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_772 = 8'h4 == inBytes_3 ? 8'hf2 : _GEN_771; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_773 = 8'h5 == inBytes_3 ? 8'h6b : _GEN_772; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_774 = 8'h6 == inBytes_3 ? 8'h6f : _GEN_773; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_775 = 8'h7 == inBytes_3 ? 8'hc5 : _GEN_774; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_776 = 8'h8 == inBytes_3 ? 8'h30 : _GEN_775; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_777 = 8'h9 == inBytes_3 ? 8'h1 : _GEN_776; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_778 = 8'ha == inBytes_3 ? 8'h67 : _GEN_777; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_779 = 8'hb == inBytes_3 ? 8'h2b : _GEN_778; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_780 = 8'hc == inBytes_3 ? 8'hfe : _GEN_779; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_781 = 8'hd == inBytes_3 ? 8'hd7 : _GEN_780; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_782 = 8'he == inBytes_3 ? 8'hab : _GEN_781; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_783 = 8'hf == inBytes_3 ? 8'h76 : _GEN_782; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_784 = 8'h10 == inBytes_3 ? 8'hca : _GEN_783; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_785 = 8'h11 == inBytes_3 ? 8'h82 : _GEN_784; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_786 = 8'h12 == inBytes_3 ? 8'hc9 : _GEN_785; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_787 = 8'h13 == inBytes_3 ? 8'h7d : _GEN_786; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_788 = 8'h14 == inBytes_3 ? 8'hfa : _GEN_787; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_789 = 8'h15 == inBytes_3 ? 8'h59 : _GEN_788; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_790 = 8'h16 == inBytes_3 ? 8'h47 : _GEN_789; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_791 = 8'h17 == inBytes_3 ? 8'hf0 : _GEN_790; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_792 = 8'h18 == inBytes_3 ? 8'had : _GEN_791; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_793 = 8'h19 == inBytes_3 ? 8'hd4 : _GEN_792; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_794 = 8'h1a == inBytes_3 ? 8'ha2 : _GEN_793; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_795 = 8'h1b == inBytes_3 ? 8'haf : _GEN_794; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_796 = 8'h1c == inBytes_3 ? 8'h9c : _GEN_795; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_797 = 8'h1d == inBytes_3 ? 8'ha4 : _GEN_796; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_798 = 8'h1e == inBytes_3 ? 8'h72 : _GEN_797; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_799 = 8'h1f == inBytes_3 ? 8'hc0 : _GEN_798; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_800 = 8'h20 == inBytes_3 ? 8'hb7 : _GEN_799; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_801 = 8'h21 == inBytes_3 ? 8'hfd : _GEN_800; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_802 = 8'h22 == inBytes_3 ? 8'h93 : _GEN_801; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_803 = 8'h23 == inBytes_3 ? 8'h26 : _GEN_802; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_804 = 8'h24 == inBytes_3 ? 8'h36 : _GEN_803; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_805 = 8'h25 == inBytes_3 ? 8'h3f : _GEN_804; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_806 = 8'h26 == inBytes_3 ? 8'hf7 : _GEN_805; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_807 = 8'h27 == inBytes_3 ? 8'hcc : _GEN_806; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_808 = 8'h28 == inBytes_3 ? 8'h34 : _GEN_807; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_809 = 8'h29 == inBytes_3 ? 8'ha5 : _GEN_808; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_810 = 8'h2a == inBytes_3 ? 8'he5 : _GEN_809; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_811 = 8'h2b == inBytes_3 ? 8'hf1 : _GEN_810; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_812 = 8'h2c == inBytes_3 ? 8'h71 : _GEN_811; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_813 = 8'h2d == inBytes_3 ? 8'hd8 : _GEN_812; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_814 = 8'h2e == inBytes_3 ? 8'h31 : _GEN_813; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_815 = 8'h2f == inBytes_3 ? 8'h15 : _GEN_814; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_816 = 8'h30 == inBytes_3 ? 8'h4 : _GEN_815; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_817 = 8'h31 == inBytes_3 ? 8'hc7 : _GEN_816; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_818 = 8'h32 == inBytes_3 ? 8'h23 : _GEN_817; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_819 = 8'h33 == inBytes_3 ? 8'hc3 : _GEN_818; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_820 = 8'h34 == inBytes_3 ? 8'h18 : _GEN_819; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_821 = 8'h35 == inBytes_3 ? 8'h96 : _GEN_820; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_822 = 8'h36 == inBytes_3 ? 8'h5 : _GEN_821; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_823 = 8'h37 == inBytes_3 ? 8'h9a : _GEN_822; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_824 = 8'h38 == inBytes_3 ? 8'h7 : _GEN_823; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_825 = 8'h39 == inBytes_3 ? 8'h12 : _GEN_824; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_826 = 8'h3a == inBytes_3 ? 8'h80 : _GEN_825; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_827 = 8'h3b == inBytes_3 ? 8'he2 : _GEN_826; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_828 = 8'h3c == inBytes_3 ? 8'heb : _GEN_827; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_829 = 8'h3d == inBytes_3 ? 8'h27 : _GEN_828; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_830 = 8'h3e == inBytes_3 ? 8'hb2 : _GEN_829; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_831 = 8'h3f == inBytes_3 ? 8'h75 : _GEN_830; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_832 = 8'h40 == inBytes_3 ? 8'h9 : _GEN_831; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_833 = 8'h41 == inBytes_3 ? 8'h83 : _GEN_832; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_834 = 8'h42 == inBytes_3 ? 8'h2c : _GEN_833; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_835 = 8'h43 == inBytes_3 ? 8'h1a : _GEN_834; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_836 = 8'h44 == inBytes_3 ? 8'h1b : _GEN_835; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_837 = 8'h45 == inBytes_3 ? 8'h6e : _GEN_836; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_838 = 8'h46 == inBytes_3 ? 8'h5a : _GEN_837; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_839 = 8'h47 == inBytes_3 ? 8'ha0 : _GEN_838; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_840 = 8'h48 == inBytes_3 ? 8'h52 : _GEN_839; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_841 = 8'h49 == inBytes_3 ? 8'h3b : _GEN_840; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_842 = 8'h4a == inBytes_3 ? 8'hd6 : _GEN_841; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_843 = 8'h4b == inBytes_3 ? 8'hb3 : _GEN_842; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_844 = 8'h4c == inBytes_3 ? 8'h29 : _GEN_843; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_845 = 8'h4d == inBytes_3 ? 8'he3 : _GEN_844; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_846 = 8'h4e == inBytes_3 ? 8'h2f : _GEN_845; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_847 = 8'h4f == inBytes_3 ? 8'h84 : _GEN_846; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_848 = 8'h50 == inBytes_3 ? 8'h53 : _GEN_847; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_849 = 8'h51 == inBytes_3 ? 8'hd1 : _GEN_848; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_850 = 8'h52 == inBytes_3 ? 8'h0 : _GEN_849; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_851 = 8'h53 == inBytes_3 ? 8'hed : _GEN_850; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_852 = 8'h54 == inBytes_3 ? 8'h20 : _GEN_851; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_853 = 8'h55 == inBytes_3 ? 8'hfc : _GEN_852; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_854 = 8'h56 == inBytes_3 ? 8'hb1 : _GEN_853; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_855 = 8'h57 == inBytes_3 ? 8'h5b : _GEN_854; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_856 = 8'h58 == inBytes_3 ? 8'h6a : _GEN_855; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_857 = 8'h59 == inBytes_3 ? 8'hcb : _GEN_856; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_858 = 8'h5a == inBytes_3 ? 8'hbe : _GEN_857; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_859 = 8'h5b == inBytes_3 ? 8'h39 : _GEN_858; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_860 = 8'h5c == inBytes_3 ? 8'h4a : _GEN_859; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_861 = 8'h5d == inBytes_3 ? 8'h4c : _GEN_860; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_862 = 8'h5e == inBytes_3 ? 8'h58 : _GEN_861; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_863 = 8'h5f == inBytes_3 ? 8'hcf : _GEN_862; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_864 = 8'h60 == inBytes_3 ? 8'hd0 : _GEN_863; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_865 = 8'h61 == inBytes_3 ? 8'hef : _GEN_864; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_866 = 8'h62 == inBytes_3 ? 8'haa : _GEN_865; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_867 = 8'h63 == inBytes_3 ? 8'hfb : _GEN_866; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_868 = 8'h64 == inBytes_3 ? 8'h43 : _GEN_867; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_869 = 8'h65 == inBytes_3 ? 8'h4d : _GEN_868; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_870 = 8'h66 == inBytes_3 ? 8'h33 : _GEN_869; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_871 = 8'h67 == inBytes_3 ? 8'h85 : _GEN_870; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_872 = 8'h68 == inBytes_3 ? 8'h45 : _GEN_871; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_873 = 8'h69 == inBytes_3 ? 8'hf9 : _GEN_872; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_874 = 8'h6a == inBytes_3 ? 8'h2 : _GEN_873; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_875 = 8'h6b == inBytes_3 ? 8'h7f : _GEN_874; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_876 = 8'h6c == inBytes_3 ? 8'h50 : _GEN_875; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_877 = 8'h6d == inBytes_3 ? 8'h3c : _GEN_876; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_878 = 8'h6e == inBytes_3 ? 8'h9f : _GEN_877; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_879 = 8'h6f == inBytes_3 ? 8'ha8 : _GEN_878; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_880 = 8'h70 == inBytes_3 ? 8'h51 : _GEN_879; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_881 = 8'h71 == inBytes_3 ? 8'ha3 : _GEN_880; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_882 = 8'h72 == inBytes_3 ? 8'h40 : _GEN_881; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_883 = 8'h73 == inBytes_3 ? 8'h8f : _GEN_882; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_884 = 8'h74 == inBytes_3 ? 8'h92 : _GEN_883; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_885 = 8'h75 == inBytes_3 ? 8'h9d : _GEN_884; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_886 = 8'h76 == inBytes_3 ? 8'h38 : _GEN_885; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_887 = 8'h77 == inBytes_3 ? 8'hf5 : _GEN_886; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_888 = 8'h78 == inBytes_3 ? 8'hbc : _GEN_887; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_889 = 8'h79 == inBytes_3 ? 8'hb6 : _GEN_888; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_890 = 8'h7a == inBytes_3 ? 8'hda : _GEN_889; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_891 = 8'h7b == inBytes_3 ? 8'h21 : _GEN_890; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_892 = 8'h7c == inBytes_3 ? 8'h10 : _GEN_891; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_893 = 8'h7d == inBytes_3 ? 8'hff : _GEN_892; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_894 = 8'h7e == inBytes_3 ? 8'hf3 : _GEN_893; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_895 = 8'h7f == inBytes_3 ? 8'hd2 : _GEN_894; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_896 = 8'h80 == inBytes_3 ? 8'hcd : _GEN_895; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_897 = 8'h81 == inBytes_3 ? 8'hc : _GEN_896; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_898 = 8'h82 == inBytes_3 ? 8'h13 : _GEN_897; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_899 = 8'h83 == inBytes_3 ? 8'hec : _GEN_898; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_900 = 8'h84 == inBytes_3 ? 8'h5f : _GEN_899; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_901 = 8'h85 == inBytes_3 ? 8'h97 : _GEN_900; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_902 = 8'h86 == inBytes_3 ? 8'h44 : _GEN_901; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_903 = 8'h87 == inBytes_3 ? 8'h17 : _GEN_902; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_904 = 8'h88 == inBytes_3 ? 8'hc4 : _GEN_903; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_905 = 8'h89 == inBytes_3 ? 8'ha7 : _GEN_904; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_906 = 8'h8a == inBytes_3 ? 8'h7e : _GEN_905; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_907 = 8'h8b == inBytes_3 ? 8'h3d : _GEN_906; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_908 = 8'h8c == inBytes_3 ? 8'h64 : _GEN_907; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_909 = 8'h8d == inBytes_3 ? 8'h5d : _GEN_908; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_910 = 8'h8e == inBytes_3 ? 8'h19 : _GEN_909; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_911 = 8'h8f == inBytes_3 ? 8'h73 : _GEN_910; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_912 = 8'h90 == inBytes_3 ? 8'h60 : _GEN_911; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_913 = 8'h91 == inBytes_3 ? 8'h81 : _GEN_912; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_914 = 8'h92 == inBytes_3 ? 8'h4f : _GEN_913; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_915 = 8'h93 == inBytes_3 ? 8'hdc : _GEN_914; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_916 = 8'h94 == inBytes_3 ? 8'h22 : _GEN_915; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_917 = 8'h95 == inBytes_3 ? 8'h2a : _GEN_916; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_918 = 8'h96 == inBytes_3 ? 8'h90 : _GEN_917; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_919 = 8'h97 == inBytes_3 ? 8'h88 : _GEN_918; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_920 = 8'h98 == inBytes_3 ? 8'h46 : _GEN_919; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_921 = 8'h99 == inBytes_3 ? 8'hee : _GEN_920; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_922 = 8'h9a == inBytes_3 ? 8'hb8 : _GEN_921; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_923 = 8'h9b == inBytes_3 ? 8'h14 : _GEN_922; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_924 = 8'h9c == inBytes_3 ? 8'hde : _GEN_923; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_925 = 8'h9d == inBytes_3 ? 8'h5e : _GEN_924; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_926 = 8'h9e == inBytes_3 ? 8'hb : _GEN_925; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_927 = 8'h9f == inBytes_3 ? 8'hdb : _GEN_926; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_928 = 8'ha0 == inBytes_3 ? 8'he0 : _GEN_927; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_929 = 8'ha1 == inBytes_3 ? 8'h32 : _GEN_928; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_930 = 8'ha2 == inBytes_3 ? 8'h3a : _GEN_929; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_931 = 8'ha3 == inBytes_3 ? 8'ha : _GEN_930; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_932 = 8'ha4 == inBytes_3 ? 8'h49 : _GEN_931; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_933 = 8'ha5 == inBytes_3 ? 8'h6 : _GEN_932; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_934 = 8'ha6 == inBytes_3 ? 8'h24 : _GEN_933; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_935 = 8'ha7 == inBytes_3 ? 8'h5c : _GEN_934; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_936 = 8'ha8 == inBytes_3 ? 8'hc2 : _GEN_935; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_937 = 8'ha9 == inBytes_3 ? 8'hd3 : _GEN_936; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_938 = 8'haa == inBytes_3 ? 8'hac : _GEN_937; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_939 = 8'hab == inBytes_3 ? 8'h62 : _GEN_938; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_940 = 8'hac == inBytes_3 ? 8'h91 : _GEN_939; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_941 = 8'had == inBytes_3 ? 8'h95 : _GEN_940; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_942 = 8'hae == inBytes_3 ? 8'he4 : _GEN_941; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_943 = 8'haf == inBytes_3 ? 8'h79 : _GEN_942; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_944 = 8'hb0 == inBytes_3 ? 8'he7 : _GEN_943; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_945 = 8'hb1 == inBytes_3 ? 8'hc8 : _GEN_944; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_946 = 8'hb2 == inBytes_3 ? 8'h37 : _GEN_945; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_947 = 8'hb3 == inBytes_3 ? 8'h6d : _GEN_946; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_948 = 8'hb4 == inBytes_3 ? 8'h8d : _GEN_947; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_949 = 8'hb5 == inBytes_3 ? 8'hd5 : _GEN_948; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_950 = 8'hb6 == inBytes_3 ? 8'h4e : _GEN_949; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_951 = 8'hb7 == inBytes_3 ? 8'ha9 : _GEN_950; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_952 = 8'hb8 == inBytes_3 ? 8'h6c : _GEN_951; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_953 = 8'hb9 == inBytes_3 ? 8'h56 : _GEN_952; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_954 = 8'hba == inBytes_3 ? 8'hf4 : _GEN_953; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_955 = 8'hbb == inBytes_3 ? 8'hea : _GEN_954; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_956 = 8'hbc == inBytes_3 ? 8'h65 : _GEN_955; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_957 = 8'hbd == inBytes_3 ? 8'h7a : _GEN_956; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_958 = 8'hbe == inBytes_3 ? 8'hae : _GEN_957; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_959 = 8'hbf == inBytes_3 ? 8'h8 : _GEN_958; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_960 = 8'hc0 == inBytes_3 ? 8'hba : _GEN_959; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_961 = 8'hc1 == inBytes_3 ? 8'h78 : _GEN_960; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_962 = 8'hc2 == inBytes_3 ? 8'h25 : _GEN_961; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_963 = 8'hc3 == inBytes_3 ? 8'h2e : _GEN_962; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_964 = 8'hc4 == inBytes_3 ? 8'h1c : _GEN_963; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_965 = 8'hc5 == inBytes_3 ? 8'ha6 : _GEN_964; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_966 = 8'hc6 == inBytes_3 ? 8'hb4 : _GEN_965; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_967 = 8'hc7 == inBytes_3 ? 8'hc6 : _GEN_966; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_968 = 8'hc8 == inBytes_3 ? 8'he8 : _GEN_967; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_969 = 8'hc9 == inBytes_3 ? 8'hdd : _GEN_968; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_970 = 8'hca == inBytes_3 ? 8'h74 : _GEN_969; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_971 = 8'hcb == inBytes_3 ? 8'h1f : _GEN_970; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_972 = 8'hcc == inBytes_3 ? 8'h4b : _GEN_971; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_973 = 8'hcd == inBytes_3 ? 8'hbd : _GEN_972; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_974 = 8'hce == inBytes_3 ? 8'h8b : _GEN_973; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_975 = 8'hcf == inBytes_3 ? 8'h8a : _GEN_974; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_976 = 8'hd0 == inBytes_3 ? 8'h70 : _GEN_975; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_977 = 8'hd1 == inBytes_3 ? 8'h3e : _GEN_976; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_978 = 8'hd2 == inBytes_3 ? 8'hb5 : _GEN_977; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_979 = 8'hd3 == inBytes_3 ? 8'h66 : _GEN_978; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_980 = 8'hd4 == inBytes_3 ? 8'h48 : _GEN_979; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_981 = 8'hd5 == inBytes_3 ? 8'h3 : _GEN_980; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_982 = 8'hd6 == inBytes_3 ? 8'hf6 : _GEN_981; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_983 = 8'hd7 == inBytes_3 ? 8'he : _GEN_982; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_984 = 8'hd8 == inBytes_3 ? 8'h61 : _GEN_983; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_985 = 8'hd9 == inBytes_3 ? 8'h35 : _GEN_984; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_986 = 8'hda == inBytes_3 ? 8'h57 : _GEN_985; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_987 = 8'hdb == inBytes_3 ? 8'hb9 : _GEN_986; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_988 = 8'hdc == inBytes_3 ? 8'h86 : _GEN_987; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_989 = 8'hdd == inBytes_3 ? 8'hc1 : _GEN_988; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_990 = 8'hde == inBytes_3 ? 8'h1d : _GEN_989; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_991 = 8'hdf == inBytes_3 ? 8'h9e : _GEN_990; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_992 = 8'he0 == inBytes_3 ? 8'he1 : _GEN_991; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_993 = 8'he1 == inBytes_3 ? 8'hf8 : _GEN_992; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_994 = 8'he2 == inBytes_3 ? 8'h98 : _GEN_993; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_995 = 8'he3 == inBytes_3 ? 8'h11 : _GEN_994; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_996 = 8'he4 == inBytes_3 ? 8'h69 : _GEN_995; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_997 = 8'he5 == inBytes_3 ? 8'hd9 : _GEN_996; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_998 = 8'he6 == inBytes_3 ? 8'h8e : _GEN_997; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_999 = 8'he7 == inBytes_3 ? 8'h94 : _GEN_998; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1000 = 8'he8 == inBytes_3 ? 8'h9b : _GEN_999; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1001 = 8'he9 == inBytes_3 ? 8'h1e : _GEN_1000; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1002 = 8'hea == inBytes_3 ? 8'h87 : _GEN_1001; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1003 = 8'heb == inBytes_3 ? 8'he9 : _GEN_1002; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1004 = 8'hec == inBytes_3 ? 8'hce : _GEN_1003; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1005 = 8'hed == inBytes_3 ? 8'h55 : _GEN_1004; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1006 = 8'hee == inBytes_3 ? 8'h28 : _GEN_1005; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1007 = 8'hef == inBytes_3 ? 8'hdf : _GEN_1006; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1008 = 8'hf0 == inBytes_3 ? 8'h8c : _GEN_1007; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1009 = 8'hf1 == inBytes_3 ? 8'ha1 : _GEN_1008; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1010 = 8'hf2 == inBytes_3 ? 8'h89 : _GEN_1009; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1011 = 8'hf3 == inBytes_3 ? 8'hd : _GEN_1010; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1012 = 8'hf4 == inBytes_3 ? 8'hbf : _GEN_1011; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1013 = 8'hf5 == inBytes_3 ? 8'he6 : _GEN_1012; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1014 = 8'hf6 == inBytes_3 ? 8'h42 : _GEN_1013; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1015 = 8'hf7 == inBytes_3 ? 8'h68 : _GEN_1014; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1016 = 8'hf8 == inBytes_3 ? 8'h41 : _GEN_1015; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1017 = 8'hf9 == inBytes_3 ? 8'h99 : _GEN_1016; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1018 = 8'hfa == inBytes_3 ? 8'h2d : _GEN_1017; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1019 = 8'hfb == inBytes_3 ? 8'hf : _GEN_1018; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1020 = 8'hfc == inBytes_3 ? 8'hb0 : _GEN_1019; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1021 = 8'hfd == inBytes_3 ? 8'h54 : _GEN_1020; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1022 = 8'hfe == inBytes_3 ? 8'hbb : _GEN_1021; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] outBytes_3 = 8'hff == inBytes_3 ? 8'h16 : _GEN_1022; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1025 = 8'h1 == inBytes_4 ? 8'h7c : 8'h63; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1026 = 8'h2 == inBytes_4 ? 8'h77 : _GEN_1025; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1027 = 8'h3 == inBytes_4 ? 8'h7b : _GEN_1026; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1028 = 8'h4 == inBytes_4 ? 8'hf2 : _GEN_1027; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1029 = 8'h5 == inBytes_4 ? 8'h6b : _GEN_1028; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1030 = 8'h6 == inBytes_4 ? 8'h6f : _GEN_1029; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1031 = 8'h7 == inBytes_4 ? 8'hc5 : _GEN_1030; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1032 = 8'h8 == inBytes_4 ? 8'h30 : _GEN_1031; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1033 = 8'h9 == inBytes_4 ? 8'h1 : _GEN_1032; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1034 = 8'ha == inBytes_4 ? 8'h67 : _GEN_1033; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1035 = 8'hb == inBytes_4 ? 8'h2b : _GEN_1034; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1036 = 8'hc == inBytes_4 ? 8'hfe : _GEN_1035; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1037 = 8'hd == inBytes_4 ? 8'hd7 : _GEN_1036; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1038 = 8'he == inBytes_4 ? 8'hab : _GEN_1037; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1039 = 8'hf == inBytes_4 ? 8'h76 : _GEN_1038; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1040 = 8'h10 == inBytes_4 ? 8'hca : _GEN_1039; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1041 = 8'h11 == inBytes_4 ? 8'h82 : _GEN_1040; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1042 = 8'h12 == inBytes_4 ? 8'hc9 : _GEN_1041; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1043 = 8'h13 == inBytes_4 ? 8'h7d : _GEN_1042; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1044 = 8'h14 == inBytes_4 ? 8'hfa : _GEN_1043; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1045 = 8'h15 == inBytes_4 ? 8'h59 : _GEN_1044; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1046 = 8'h16 == inBytes_4 ? 8'h47 : _GEN_1045; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1047 = 8'h17 == inBytes_4 ? 8'hf0 : _GEN_1046; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1048 = 8'h18 == inBytes_4 ? 8'had : _GEN_1047; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1049 = 8'h19 == inBytes_4 ? 8'hd4 : _GEN_1048; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1050 = 8'h1a == inBytes_4 ? 8'ha2 : _GEN_1049; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1051 = 8'h1b == inBytes_4 ? 8'haf : _GEN_1050; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1052 = 8'h1c == inBytes_4 ? 8'h9c : _GEN_1051; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1053 = 8'h1d == inBytes_4 ? 8'ha4 : _GEN_1052; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1054 = 8'h1e == inBytes_4 ? 8'h72 : _GEN_1053; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1055 = 8'h1f == inBytes_4 ? 8'hc0 : _GEN_1054; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1056 = 8'h20 == inBytes_4 ? 8'hb7 : _GEN_1055; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1057 = 8'h21 == inBytes_4 ? 8'hfd : _GEN_1056; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1058 = 8'h22 == inBytes_4 ? 8'h93 : _GEN_1057; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1059 = 8'h23 == inBytes_4 ? 8'h26 : _GEN_1058; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1060 = 8'h24 == inBytes_4 ? 8'h36 : _GEN_1059; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1061 = 8'h25 == inBytes_4 ? 8'h3f : _GEN_1060; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1062 = 8'h26 == inBytes_4 ? 8'hf7 : _GEN_1061; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1063 = 8'h27 == inBytes_4 ? 8'hcc : _GEN_1062; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1064 = 8'h28 == inBytes_4 ? 8'h34 : _GEN_1063; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1065 = 8'h29 == inBytes_4 ? 8'ha5 : _GEN_1064; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1066 = 8'h2a == inBytes_4 ? 8'he5 : _GEN_1065; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1067 = 8'h2b == inBytes_4 ? 8'hf1 : _GEN_1066; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1068 = 8'h2c == inBytes_4 ? 8'h71 : _GEN_1067; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1069 = 8'h2d == inBytes_4 ? 8'hd8 : _GEN_1068; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1070 = 8'h2e == inBytes_4 ? 8'h31 : _GEN_1069; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1071 = 8'h2f == inBytes_4 ? 8'h15 : _GEN_1070; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1072 = 8'h30 == inBytes_4 ? 8'h4 : _GEN_1071; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1073 = 8'h31 == inBytes_4 ? 8'hc7 : _GEN_1072; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1074 = 8'h32 == inBytes_4 ? 8'h23 : _GEN_1073; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1075 = 8'h33 == inBytes_4 ? 8'hc3 : _GEN_1074; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1076 = 8'h34 == inBytes_4 ? 8'h18 : _GEN_1075; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1077 = 8'h35 == inBytes_4 ? 8'h96 : _GEN_1076; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1078 = 8'h36 == inBytes_4 ? 8'h5 : _GEN_1077; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1079 = 8'h37 == inBytes_4 ? 8'h9a : _GEN_1078; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1080 = 8'h38 == inBytes_4 ? 8'h7 : _GEN_1079; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1081 = 8'h39 == inBytes_4 ? 8'h12 : _GEN_1080; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1082 = 8'h3a == inBytes_4 ? 8'h80 : _GEN_1081; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1083 = 8'h3b == inBytes_4 ? 8'he2 : _GEN_1082; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1084 = 8'h3c == inBytes_4 ? 8'heb : _GEN_1083; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1085 = 8'h3d == inBytes_4 ? 8'h27 : _GEN_1084; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1086 = 8'h3e == inBytes_4 ? 8'hb2 : _GEN_1085; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1087 = 8'h3f == inBytes_4 ? 8'h75 : _GEN_1086; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1088 = 8'h40 == inBytes_4 ? 8'h9 : _GEN_1087; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1089 = 8'h41 == inBytes_4 ? 8'h83 : _GEN_1088; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1090 = 8'h42 == inBytes_4 ? 8'h2c : _GEN_1089; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1091 = 8'h43 == inBytes_4 ? 8'h1a : _GEN_1090; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1092 = 8'h44 == inBytes_4 ? 8'h1b : _GEN_1091; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1093 = 8'h45 == inBytes_4 ? 8'h6e : _GEN_1092; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1094 = 8'h46 == inBytes_4 ? 8'h5a : _GEN_1093; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1095 = 8'h47 == inBytes_4 ? 8'ha0 : _GEN_1094; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1096 = 8'h48 == inBytes_4 ? 8'h52 : _GEN_1095; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1097 = 8'h49 == inBytes_4 ? 8'h3b : _GEN_1096; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1098 = 8'h4a == inBytes_4 ? 8'hd6 : _GEN_1097; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1099 = 8'h4b == inBytes_4 ? 8'hb3 : _GEN_1098; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1100 = 8'h4c == inBytes_4 ? 8'h29 : _GEN_1099; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1101 = 8'h4d == inBytes_4 ? 8'he3 : _GEN_1100; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1102 = 8'h4e == inBytes_4 ? 8'h2f : _GEN_1101; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1103 = 8'h4f == inBytes_4 ? 8'h84 : _GEN_1102; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1104 = 8'h50 == inBytes_4 ? 8'h53 : _GEN_1103; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1105 = 8'h51 == inBytes_4 ? 8'hd1 : _GEN_1104; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1106 = 8'h52 == inBytes_4 ? 8'h0 : _GEN_1105; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1107 = 8'h53 == inBytes_4 ? 8'hed : _GEN_1106; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1108 = 8'h54 == inBytes_4 ? 8'h20 : _GEN_1107; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1109 = 8'h55 == inBytes_4 ? 8'hfc : _GEN_1108; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1110 = 8'h56 == inBytes_4 ? 8'hb1 : _GEN_1109; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1111 = 8'h57 == inBytes_4 ? 8'h5b : _GEN_1110; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1112 = 8'h58 == inBytes_4 ? 8'h6a : _GEN_1111; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1113 = 8'h59 == inBytes_4 ? 8'hcb : _GEN_1112; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1114 = 8'h5a == inBytes_4 ? 8'hbe : _GEN_1113; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1115 = 8'h5b == inBytes_4 ? 8'h39 : _GEN_1114; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1116 = 8'h5c == inBytes_4 ? 8'h4a : _GEN_1115; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1117 = 8'h5d == inBytes_4 ? 8'h4c : _GEN_1116; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1118 = 8'h5e == inBytes_4 ? 8'h58 : _GEN_1117; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1119 = 8'h5f == inBytes_4 ? 8'hcf : _GEN_1118; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1120 = 8'h60 == inBytes_4 ? 8'hd0 : _GEN_1119; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1121 = 8'h61 == inBytes_4 ? 8'hef : _GEN_1120; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1122 = 8'h62 == inBytes_4 ? 8'haa : _GEN_1121; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1123 = 8'h63 == inBytes_4 ? 8'hfb : _GEN_1122; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1124 = 8'h64 == inBytes_4 ? 8'h43 : _GEN_1123; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1125 = 8'h65 == inBytes_4 ? 8'h4d : _GEN_1124; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1126 = 8'h66 == inBytes_4 ? 8'h33 : _GEN_1125; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1127 = 8'h67 == inBytes_4 ? 8'h85 : _GEN_1126; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1128 = 8'h68 == inBytes_4 ? 8'h45 : _GEN_1127; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1129 = 8'h69 == inBytes_4 ? 8'hf9 : _GEN_1128; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1130 = 8'h6a == inBytes_4 ? 8'h2 : _GEN_1129; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1131 = 8'h6b == inBytes_4 ? 8'h7f : _GEN_1130; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1132 = 8'h6c == inBytes_4 ? 8'h50 : _GEN_1131; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1133 = 8'h6d == inBytes_4 ? 8'h3c : _GEN_1132; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1134 = 8'h6e == inBytes_4 ? 8'h9f : _GEN_1133; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1135 = 8'h6f == inBytes_4 ? 8'ha8 : _GEN_1134; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1136 = 8'h70 == inBytes_4 ? 8'h51 : _GEN_1135; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1137 = 8'h71 == inBytes_4 ? 8'ha3 : _GEN_1136; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1138 = 8'h72 == inBytes_4 ? 8'h40 : _GEN_1137; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1139 = 8'h73 == inBytes_4 ? 8'h8f : _GEN_1138; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1140 = 8'h74 == inBytes_4 ? 8'h92 : _GEN_1139; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1141 = 8'h75 == inBytes_4 ? 8'h9d : _GEN_1140; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1142 = 8'h76 == inBytes_4 ? 8'h38 : _GEN_1141; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1143 = 8'h77 == inBytes_4 ? 8'hf5 : _GEN_1142; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1144 = 8'h78 == inBytes_4 ? 8'hbc : _GEN_1143; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1145 = 8'h79 == inBytes_4 ? 8'hb6 : _GEN_1144; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1146 = 8'h7a == inBytes_4 ? 8'hda : _GEN_1145; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1147 = 8'h7b == inBytes_4 ? 8'h21 : _GEN_1146; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1148 = 8'h7c == inBytes_4 ? 8'h10 : _GEN_1147; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1149 = 8'h7d == inBytes_4 ? 8'hff : _GEN_1148; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1150 = 8'h7e == inBytes_4 ? 8'hf3 : _GEN_1149; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1151 = 8'h7f == inBytes_4 ? 8'hd2 : _GEN_1150; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1152 = 8'h80 == inBytes_4 ? 8'hcd : _GEN_1151; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1153 = 8'h81 == inBytes_4 ? 8'hc : _GEN_1152; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1154 = 8'h82 == inBytes_4 ? 8'h13 : _GEN_1153; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1155 = 8'h83 == inBytes_4 ? 8'hec : _GEN_1154; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1156 = 8'h84 == inBytes_4 ? 8'h5f : _GEN_1155; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1157 = 8'h85 == inBytes_4 ? 8'h97 : _GEN_1156; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1158 = 8'h86 == inBytes_4 ? 8'h44 : _GEN_1157; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1159 = 8'h87 == inBytes_4 ? 8'h17 : _GEN_1158; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1160 = 8'h88 == inBytes_4 ? 8'hc4 : _GEN_1159; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1161 = 8'h89 == inBytes_4 ? 8'ha7 : _GEN_1160; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1162 = 8'h8a == inBytes_4 ? 8'h7e : _GEN_1161; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1163 = 8'h8b == inBytes_4 ? 8'h3d : _GEN_1162; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1164 = 8'h8c == inBytes_4 ? 8'h64 : _GEN_1163; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1165 = 8'h8d == inBytes_4 ? 8'h5d : _GEN_1164; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1166 = 8'h8e == inBytes_4 ? 8'h19 : _GEN_1165; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1167 = 8'h8f == inBytes_4 ? 8'h73 : _GEN_1166; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1168 = 8'h90 == inBytes_4 ? 8'h60 : _GEN_1167; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1169 = 8'h91 == inBytes_4 ? 8'h81 : _GEN_1168; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1170 = 8'h92 == inBytes_4 ? 8'h4f : _GEN_1169; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1171 = 8'h93 == inBytes_4 ? 8'hdc : _GEN_1170; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1172 = 8'h94 == inBytes_4 ? 8'h22 : _GEN_1171; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1173 = 8'h95 == inBytes_4 ? 8'h2a : _GEN_1172; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1174 = 8'h96 == inBytes_4 ? 8'h90 : _GEN_1173; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1175 = 8'h97 == inBytes_4 ? 8'h88 : _GEN_1174; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1176 = 8'h98 == inBytes_4 ? 8'h46 : _GEN_1175; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1177 = 8'h99 == inBytes_4 ? 8'hee : _GEN_1176; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1178 = 8'h9a == inBytes_4 ? 8'hb8 : _GEN_1177; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1179 = 8'h9b == inBytes_4 ? 8'h14 : _GEN_1178; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1180 = 8'h9c == inBytes_4 ? 8'hde : _GEN_1179; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1181 = 8'h9d == inBytes_4 ? 8'h5e : _GEN_1180; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1182 = 8'h9e == inBytes_4 ? 8'hb : _GEN_1181; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1183 = 8'h9f == inBytes_4 ? 8'hdb : _GEN_1182; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1184 = 8'ha0 == inBytes_4 ? 8'he0 : _GEN_1183; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1185 = 8'ha1 == inBytes_4 ? 8'h32 : _GEN_1184; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1186 = 8'ha2 == inBytes_4 ? 8'h3a : _GEN_1185; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1187 = 8'ha3 == inBytes_4 ? 8'ha : _GEN_1186; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1188 = 8'ha4 == inBytes_4 ? 8'h49 : _GEN_1187; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1189 = 8'ha5 == inBytes_4 ? 8'h6 : _GEN_1188; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1190 = 8'ha6 == inBytes_4 ? 8'h24 : _GEN_1189; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1191 = 8'ha7 == inBytes_4 ? 8'h5c : _GEN_1190; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1192 = 8'ha8 == inBytes_4 ? 8'hc2 : _GEN_1191; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1193 = 8'ha9 == inBytes_4 ? 8'hd3 : _GEN_1192; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1194 = 8'haa == inBytes_4 ? 8'hac : _GEN_1193; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1195 = 8'hab == inBytes_4 ? 8'h62 : _GEN_1194; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1196 = 8'hac == inBytes_4 ? 8'h91 : _GEN_1195; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1197 = 8'had == inBytes_4 ? 8'h95 : _GEN_1196; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1198 = 8'hae == inBytes_4 ? 8'he4 : _GEN_1197; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1199 = 8'haf == inBytes_4 ? 8'h79 : _GEN_1198; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1200 = 8'hb0 == inBytes_4 ? 8'he7 : _GEN_1199; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1201 = 8'hb1 == inBytes_4 ? 8'hc8 : _GEN_1200; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1202 = 8'hb2 == inBytes_4 ? 8'h37 : _GEN_1201; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1203 = 8'hb3 == inBytes_4 ? 8'h6d : _GEN_1202; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1204 = 8'hb4 == inBytes_4 ? 8'h8d : _GEN_1203; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1205 = 8'hb5 == inBytes_4 ? 8'hd5 : _GEN_1204; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1206 = 8'hb6 == inBytes_4 ? 8'h4e : _GEN_1205; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1207 = 8'hb7 == inBytes_4 ? 8'ha9 : _GEN_1206; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1208 = 8'hb8 == inBytes_4 ? 8'h6c : _GEN_1207; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1209 = 8'hb9 == inBytes_4 ? 8'h56 : _GEN_1208; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1210 = 8'hba == inBytes_4 ? 8'hf4 : _GEN_1209; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1211 = 8'hbb == inBytes_4 ? 8'hea : _GEN_1210; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1212 = 8'hbc == inBytes_4 ? 8'h65 : _GEN_1211; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1213 = 8'hbd == inBytes_4 ? 8'h7a : _GEN_1212; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1214 = 8'hbe == inBytes_4 ? 8'hae : _GEN_1213; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1215 = 8'hbf == inBytes_4 ? 8'h8 : _GEN_1214; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1216 = 8'hc0 == inBytes_4 ? 8'hba : _GEN_1215; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1217 = 8'hc1 == inBytes_4 ? 8'h78 : _GEN_1216; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1218 = 8'hc2 == inBytes_4 ? 8'h25 : _GEN_1217; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1219 = 8'hc3 == inBytes_4 ? 8'h2e : _GEN_1218; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1220 = 8'hc4 == inBytes_4 ? 8'h1c : _GEN_1219; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1221 = 8'hc5 == inBytes_4 ? 8'ha6 : _GEN_1220; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1222 = 8'hc6 == inBytes_4 ? 8'hb4 : _GEN_1221; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1223 = 8'hc7 == inBytes_4 ? 8'hc6 : _GEN_1222; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1224 = 8'hc8 == inBytes_4 ? 8'he8 : _GEN_1223; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1225 = 8'hc9 == inBytes_4 ? 8'hdd : _GEN_1224; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1226 = 8'hca == inBytes_4 ? 8'h74 : _GEN_1225; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1227 = 8'hcb == inBytes_4 ? 8'h1f : _GEN_1226; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1228 = 8'hcc == inBytes_4 ? 8'h4b : _GEN_1227; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1229 = 8'hcd == inBytes_4 ? 8'hbd : _GEN_1228; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1230 = 8'hce == inBytes_4 ? 8'h8b : _GEN_1229; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1231 = 8'hcf == inBytes_4 ? 8'h8a : _GEN_1230; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1232 = 8'hd0 == inBytes_4 ? 8'h70 : _GEN_1231; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1233 = 8'hd1 == inBytes_4 ? 8'h3e : _GEN_1232; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1234 = 8'hd2 == inBytes_4 ? 8'hb5 : _GEN_1233; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1235 = 8'hd3 == inBytes_4 ? 8'h66 : _GEN_1234; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1236 = 8'hd4 == inBytes_4 ? 8'h48 : _GEN_1235; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1237 = 8'hd5 == inBytes_4 ? 8'h3 : _GEN_1236; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1238 = 8'hd6 == inBytes_4 ? 8'hf6 : _GEN_1237; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1239 = 8'hd7 == inBytes_4 ? 8'he : _GEN_1238; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1240 = 8'hd8 == inBytes_4 ? 8'h61 : _GEN_1239; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1241 = 8'hd9 == inBytes_4 ? 8'h35 : _GEN_1240; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1242 = 8'hda == inBytes_4 ? 8'h57 : _GEN_1241; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1243 = 8'hdb == inBytes_4 ? 8'hb9 : _GEN_1242; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1244 = 8'hdc == inBytes_4 ? 8'h86 : _GEN_1243; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1245 = 8'hdd == inBytes_4 ? 8'hc1 : _GEN_1244; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1246 = 8'hde == inBytes_4 ? 8'h1d : _GEN_1245; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1247 = 8'hdf == inBytes_4 ? 8'h9e : _GEN_1246; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1248 = 8'he0 == inBytes_4 ? 8'he1 : _GEN_1247; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1249 = 8'he1 == inBytes_4 ? 8'hf8 : _GEN_1248; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1250 = 8'he2 == inBytes_4 ? 8'h98 : _GEN_1249; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1251 = 8'he3 == inBytes_4 ? 8'h11 : _GEN_1250; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1252 = 8'he4 == inBytes_4 ? 8'h69 : _GEN_1251; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1253 = 8'he5 == inBytes_4 ? 8'hd9 : _GEN_1252; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1254 = 8'he6 == inBytes_4 ? 8'h8e : _GEN_1253; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1255 = 8'he7 == inBytes_4 ? 8'h94 : _GEN_1254; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1256 = 8'he8 == inBytes_4 ? 8'h9b : _GEN_1255; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1257 = 8'he9 == inBytes_4 ? 8'h1e : _GEN_1256; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1258 = 8'hea == inBytes_4 ? 8'h87 : _GEN_1257; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1259 = 8'heb == inBytes_4 ? 8'he9 : _GEN_1258; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1260 = 8'hec == inBytes_4 ? 8'hce : _GEN_1259; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1261 = 8'hed == inBytes_4 ? 8'h55 : _GEN_1260; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1262 = 8'hee == inBytes_4 ? 8'h28 : _GEN_1261; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1263 = 8'hef == inBytes_4 ? 8'hdf : _GEN_1262; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1264 = 8'hf0 == inBytes_4 ? 8'h8c : _GEN_1263; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1265 = 8'hf1 == inBytes_4 ? 8'ha1 : _GEN_1264; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1266 = 8'hf2 == inBytes_4 ? 8'h89 : _GEN_1265; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1267 = 8'hf3 == inBytes_4 ? 8'hd : _GEN_1266; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1268 = 8'hf4 == inBytes_4 ? 8'hbf : _GEN_1267; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1269 = 8'hf5 == inBytes_4 ? 8'he6 : _GEN_1268; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1270 = 8'hf6 == inBytes_4 ? 8'h42 : _GEN_1269; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1271 = 8'hf7 == inBytes_4 ? 8'h68 : _GEN_1270; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1272 = 8'hf8 == inBytes_4 ? 8'h41 : _GEN_1271; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1273 = 8'hf9 == inBytes_4 ? 8'h99 : _GEN_1272; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1274 = 8'hfa == inBytes_4 ? 8'h2d : _GEN_1273; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1275 = 8'hfb == inBytes_4 ? 8'hf : _GEN_1274; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1276 = 8'hfc == inBytes_4 ? 8'hb0 : _GEN_1275; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1277 = 8'hfd == inBytes_4 ? 8'h54 : _GEN_1276; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1278 = 8'hfe == inBytes_4 ? 8'hbb : _GEN_1277; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] outBytes_4 = 8'hff == inBytes_4 ? 8'h16 : _GEN_1278; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1281 = 8'h1 == inBytes_5 ? 8'h7c : 8'h63; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1282 = 8'h2 == inBytes_5 ? 8'h77 : _GEN_1281; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1283 = 8'h3 == inBytes_5 ? 8'h7b : _GEN_1282; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1284 = 8'h4 == inBytes_5 ? 8'hf2 : _GEN_1283; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1285 = 8'h5 == inBytes_5 ? 8'h6b : _GEN_1284; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1286 = 8'h6 == inBytes_5 ? 8'h6f : _GEN_1285; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1287 = 8'h7 == inBytes_5 ? 8'hc5 : _GEN_1286; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1288 = 8'h8 == inBytes_5 ? 8'h30 : _GEN_1287; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1289 = 8'h9 == inBytes_5 ? 8'h1 : _GEN_1288; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1290 = 8'ha == inBytes_5 ? 8'h67 : _GEN_1289; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1291 = 8'hb == inBytes_5 ? 8'h2b : _GEN_1290; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1292 = 8'hc == inBytes_5 ? 8'hfe : _GEN_1291; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1293 = 8'hd == inBytes_5 ? 8'hd7 : _GEN_1292; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1294 = 8'he == inBytes_5 ? 8'hab : _GEN_1293; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1295 = 8'hf == inBytes_5 ? 8'h76 : _GEN_1294; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1296 = 8'h10 == inBytes_5 ? 8'hca : _GEN_1295; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1297 = 8'h11 == inBytes_5 ? 8'h82 : _GEN_1296; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1298 = 8'h12 == inBytes_5 ? 8'hc9 : _GEN_1297; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1299 = 8'h13 == inBytes_5 ? 8'h7d : _GEN_1298; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1300 = 8'h14 == inBytes_5 ? 8'hfa : _GEN_1299; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1301 = 8'h15 == inBytes_5 ? 8'h59 : _GEN_1300; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1302 = 8'h16 == inBytes_5 ? 8'h47 : _GEN_1301; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1303 = 8'h17 == inBytes_5 ? 8'hf0 : _GEN_1302; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1304 = 8'h18 == inBytes_5 ? 8'had : _GEN_1303; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1305 = 8'h19 == inBytes_5 ? 8'hd4 : _GEN_1304; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1306 = 8'h1a == inBytes_5 ? 8'ha2 : _GEN_1305; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1307 = 8'h1b == inBytes_5 ? 8'haf : _GEN_1306; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1308 = 8'h1c == inBytes_5 ? 8'h9c : _GEN_1307; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1309 = 8'h1d == inBytes_5 ? 8'ha4 : _GEN_1308; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1310 = 8'h1e == inBytes_5 ? 8'h72 : _GEN_1309; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1311 = 8'h1f == inBytes_5 ? 8'hc0 : _GEN_1310; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1312 = 8'h20 == inBytes_5 ? 8'hb7 : _GEN_1311; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1313 = 8'h21 == inBytes_5 ? 8'hfd : _GEN_1312; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1314 = 8'h22 == inBytes_5 ? 8'h93 : _GEN_1313; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1315 = 8'h23 == inBytes_5 ? 8'h26 : _GEN_1314; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1316 = 8'h24 == inBytes_5 ? 8'h36 : _GEN_1315; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1317 = 8'h25 == inBytes_5 ? 8'h3f : _GEN_1316; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1318 = 8'h26 == inBytes_5 ? 8'hf7 : _GEN_1317; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1319 = 8'h27 == inBytes_5 ? 8'hcc : _GEN_1318; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1320 = 8'h28 == inBytes_5 ? 8'h34 : _GEN_1319; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1321 = 8'h29 == inBytes_5 ? 8'ha5 : _GEN_1320; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1322 = 8'h2a == inBytes_5 ? 8'he5 : _GEN_1321; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1323 = 8'h2b == inBytes_5 ? 8'hf1 : _GEN_1322; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1324 = 8'h2c == inBytes_5 ? 8'h71 : _GEN_1323; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1325 = 8'h2d == inBytes_5 ? 8'hd8 : _GEN_1324; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1326 = 8'h2e == inBytes_5 ? 8'h31 : _GEN_1325; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1327 = 8'h2f == inBytes_5 ? 8'h15 : _GEN_1326; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1328 = 8'h30 == inBytes_5 ? 8'h4 : _GEN_1327; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1329 = 8'h31 == inBytes_5 ? 8'hc7 : _GEN_1328; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1330 = 8'h32 == inBytes_5 ? 8'h23 : _GEN_1329; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1331 = 8'h33 == inBytes_5 ? 8'hc3 : _GEN_1330; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1332 = 8'h34 == inBytes_5 ? 8'h18 : _GEN_1331; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1333 = 8'h35 == inBytes_5 ? 8'h96 : _GEN_1332; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1334 = 8'h36 == inBytes_5 ? 8'h5 : _GEN_1333; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1335 = 8'h37 == inBytes_5 ? 8'h9a : _GEN_1334; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1336 = 8'h38 == inBytes_5 ? 8'h7 : _GEN_1335; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1337 = 8'h39 == inBytes_5 ? 8'h12 : _GEN_1336; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1338 = 8'h3a == inBytes_5 ? 8'h80 : _GEN_1337; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1339 = 8'h3b == inBytes_5 ? 8'he2 : _GEN_1338; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1340 = 8'h3c == inBytes_5 ? 8'heb : _GEN_1339; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1341 = 8'h3d == inBytes_5 ? 8'h27 : _GEN_1340; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1342 = 8'h3e == inBytes_5 ? 8'hb2 : _GEN_1341; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1343 = 8'h3f == inBytes_5 ? 8'h75 : _GEN_1342; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1344 = 8'h40 == inBytes_5 ? 8'h9 : _GEN_1343; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1345 = 8'h41 == inBytes_5 ? 8'h83 : _GEN_1344; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1346 = 8'h42 == inBytes_5 ? 8'h2c : _GEN_1345; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1347 = 8'h43 == inBytes_5 ? 8'h1a : _GEN_1346; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1348 = 8'h44 == inBytes_5 ? 8'h1b : _GEN_1347; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1349 = 8'h45 == inBytes_5 ? 8'h6e : _GEN_1348; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1350 = 8'h46 == inBytes_5 ? 8'h5a : _GEN_1349; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1351 = 8'h47 == inBytes_5 ? 8'ha0 : _GEN_1350; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1352 = 8'h48 == inBytes_5 ? 8'h52 : _GEN_1351; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1353 = 8'h49 == inBytes_5 ? 8'h3b : _GEN_1352; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1354 = 8'h4a == inBytes_5 ? 8'hd6 : _GEN_1353; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1355 = 8'h4b == inBytes_5 ? 8'hb3 : _GEN_1354; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1356 = 8'h4c == inBytes_5 ? 8'h29 : _GEN_1355; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1357 = 8'h4d == inBytes_5 ? 8'he3 : _GEN_1356; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1358 = 8'h4e == inBytes_5 ? 8'h2f : _GEN_1357; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1359 = 8'h4f == inBytes_5 ? 8'h84 : _GEN_1358; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1360 = 8'h50 == inBytes_5 ? 8'h53 : _GEN_1359; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1361 = 8'h51 == inBytes_5 ? 8'hd1 : _GEN_1360; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1362 = 8'h52 == inBytes_5 ? 8'h0 : _GEN_1361; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1363 = 8'h53 == inBytes_5 ? 8'hed : _GEN_1362; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1364 = 8'h54 == inBytes_5 ? 8'h20 : _GEN_1363; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1365 = 8'h55 == inBytes_5 ? 8'hfc : _GEN_1364; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1366 = 8'h56 == inBytes_5 ? 8'hb1 : _GEN_1365; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1367 = 8'h57 == inBytes_5 ? 8'h5b : _GEN_1366; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1368 = 8'h58 == inBytes_5 ? 8'h6a : _GEN_1367; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1369 = 8'h59 == inBytes_5 ? 8'hcb : _GEN_1368; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1370 = 8'h5a == inBytes_5 ? 8'hbe : _GEN_1369; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1371 = 8'h5b == inBytes_5 ? 8'h39 : _GEN_1370; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1372 = 8'h5c == inBytes_5 ? 8'h4a : _GEN_1371; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1373 = 8'h5d == inBytes_5 ? 8'h4c : _GEN_1372; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1374 = 8'h5e == inBytes_5 ? 8'h58 : _GEN_1373; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1375 = 8'h5f == inBytes_5 ? 8'hcf : _GEN_1374; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1376 = 8'h60 == inBytes_5 ? 8'hd0 : _GEN_1375; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1377 = 8'h61 == inBytes_5 ? 8'hef : _GEN_1376; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1378 = 8'h62 == inBytes_5 ? 8'haa : _GEN_1377; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1379 = 8'h63 == inBytes_5 ? 8'hfb : _GEN_1378; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1380 = 8'h64 == inBytes_5 ? 8'h43 : _GEN_1379; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1381 = 8'h65 == inBytes_5 ? 8'h4d : _GEN_1380; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1382 = 8'h66 == inBytes_5 ? 8'h33 : _GEN_1381; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1383 = 8'h67 == inBytes_5 ? 8'h85 : _GEN_1382; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1384 = 8'h68 == inBytes_5 ? 8'h45 : _GEN_1383; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1385 = 8'h69 == inBytes_5 ? 8'hf9 : _GEN_1384; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1386 = 8'h6a == inBytes_5 ? 8'h2 : _GEN_1385; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1387 = 8'h6b == inBytes_5 ? 8'h7f : _GEN_1386; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1388 = 8'h6c == inBytes_5 ? 8'h50 : _GEN_1387; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1389 = 8'h6d == inBytes_5 ? 8'h3c : _GEN_1388; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1390 = 8'h6e == inBytes_5 ? 8'h9f : _GEN_1389; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1391 = 8'h6f == inBytes_5 ? 8'ha8 : _GEN_1390; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1392 = 8'h70 == inBytes_5 ? 8'h51 : _GEN_1391; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1393 = 8'h71 == inBytes_5 ? 8'ha3 : _GEN_1392; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1394 = 8'h72 == inBytes_5 ? 8'h40 : _GEN_1393; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1395 = 8'h73 == inBytes_5 ? 8'h8f : _GEN_1394; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1396 = 8'h74 == inBytes_5 ? 8'h92 : _GEN_1395; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1397 = 8'h75 == inBytes_5 ? 8'h9d : _GEN_1396; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1398 = 8'h76 == inBytes_5 ? 8'h38 : _GEN_1397; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1399 = 8'h77 == inBytes_5 ? 8'hf5 : _GEN_1398; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1400 = 8'h78 == inBytes_5 ? 8'hbc : _GEN_1399; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1401 = 8'h79 == inBytes_5 ? 8'hb6 : _GEN_1400; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1402 = 8'h7a == inBytes_5 ? 8'hda : _GEN_1401; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1403 = 8'h7b == inBytes_5 ? 8'h21 : _GEN_1402; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1404 = 8'h7c == inBytes_5 ? 8'h10 : _GEN_1403; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1405 = 8'h7d == inBytes_5 ? 8'hff : _GEN_1404; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1406 = 8'h7e == inBytes_5 ? 8'hf3 : _GEN_1405; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1407 = 8'h7f == inBytes_5 ? 8'hd2 : _GEN_1406; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1408 = 8'h80 == inBytes_5 ? 8'hcd : _GEN_1407; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1409 = 8'h81 == inBytes_5 ? 8'hc : _GEN_1408; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1410 = 8'h82 == inBytes_5 ? 8'h13 : _GEN_1409; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1411 = 8'h83 == inBytes_5 ? 8'hec : _GEN_1410; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1412 = 8'h84 == inBytes_5 ? 8'h5f : _GEN_1411; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1413 = 8'h85 == inBytes_5 ? 8'h97 : _GEN_1412; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1414 = 8'h86 == inBytes_5 ? 8'h44 : _GEN_1413; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1415 = 8'h87 == inBytes_5 ? 8'h17 : _GEN_1414; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1416 = 8'h88 == inBytes_5 ? 8'hc4 : _GEN_1415; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1417 = 8'h89 == inBytes_5 ? 8'ha7 : _GEN_1416; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1418 = 8'h8a == inBytes_5 ? 8'h7e : _GEN_1417; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1419 = 8'h8b == inBytes_5 ? 8'h3d : _GEN_1418; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1420 = 8'h8c == inBytes_5 ? 8'h64 : _GEN_1419; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1421 = 8'h8d == inBytes_5 ? 8'h5d : _GEN_1420; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1422 = 8'h8e == inBytes_5 ? 8'h19 : _GEN_1421; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1423 = 8'h8f == inBytes_5 ? 8'h73 : _GEN_1422; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1424 = 8'h90 == inBytes_5 ? 8'h60 : _GEN_1423; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1425 = 8'h91 == inBytes_5 ? 8'h81 : _GEN_1424; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1426 = 8'h92 == inBytes_5 ? 8'h4f : _GEN_1425; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1427 = 8'h93 == inBytes_5 ? 8'hdc : _GEN_1426; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1428 = 8'h94 == inBytes_5 ? 8'h22 : _GEN_1427; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1429 = 8'h95 == inBytes_5 ? 8'h2a : _GEN_1428; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1430 = 8'h96 == inBytes_5 ? 8'h90 : _GEN_1429; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1431 = 8'h97 == inBytes_5 ? 8'h88 : _GEN_1430; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1432 = 8'h98 == inBytes_5 ? 8'h46 : _GEN_1431; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1433 = 8'h99 == inBytes_5 ? 8'hee : _GEN_1432; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1434 = 8'h9a == inBytes_5 ? 8'hb8 : _GEN_1433; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1435 = 8'h9b == inBytes_5 ? 8'h14 : _GEN_1434; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1436 = 8'h9c == inBytes_5 ? 8'hde : _GEN_1435; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1437 = 8'h9d == inBytes_5 ? 8'h5e : _GEN_1436; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1438 = 8'h9e == inBytes_5 ? 8'hb : _GEN_1437; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1439 = 8'h9f == inBytes_5 ? 8'hdb : _GEN_1438; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1440 = 8'ha0 == inBytes_5 ? 8'he0 : _GEN_1439; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1441 = 8'ha1 == inBytes_5 ? 8'h32 : _GEN_1440; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1442 = 8'ha2 == inBytes_5 ? 8'h3a : _GEN_1441; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1443 = 8'ha3 == inBytes_5 ? 8'ha : _GEN_1442; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1444 = 8'ha4 == inBytes_5 ? 8'h49 : _GEN_1443; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1445 = 8'ha5 == inBytes_5 ? 8'h6 : _GEN_1444; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1446 = 8'ha6 == inBytes_5 ? 8'h24 : _GEN_1445; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1447 = 8'ha7 == inBytes_5 ? 8'h5c : _GEN_1446; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1448 = 8'ha8 == inBytes_5 ? 8'hc2 : _GEN_1447; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1449 = 8'ha9 == inBytes_5 ? 8'hd3 : _GEN_1448; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1450 = 8'haa == inBytes_5 ? 8'hac : _GEN_1449; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1451 = 8'hab == inBytes_5 ? 8'h62 : _GEN_1450; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1452 = 8'hac == inBytes_5 ? 8'h91 : _GEN_1451; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1453 = 8'had == inBytes_5 ? 8'h95 : _GEN_1452; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1454 = 8'hae == inBytes_5 ? 8'he4 : _GEN_1453; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1455 = 8'haf == inBytes_5 ? 8'h79 : _GEN_1454; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1456 = 8'hb0 == inBytes_5 ? 8'he7 : _GEN_1455; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1457 = 8'hb1 == inBytes_5 ? 8'hc8 : _GEN_1456; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1458 = 8'hb2 == inBytes_5 ? 8'h37 : _GEN_1457; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1459 = 8'hb3 == inBytes_5 ? 8'h6d : _GEN_1458; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1460 = 8'hb4 == inBytes_5 ? 8'h8d : _GEN_1459; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1461 = 8'hb5 == inBytes_5 ? 8'hd5 : _GEN_1460; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1462 = 8'hb6 == inBytes_5 ? 8'h4e : _GEN_1461; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1463 = 8'hb7 == inBytes_5 ? 8'ha9 : _GEN_1462; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1464 = 8'hb8 == inBytes_5 ? 8'h6c : _GEN_1463; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1465 = 8'hb9 == inBytes_5 ? 8'h56 : _GEN_1464; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1466 = 8'hba == inBytes_5 ? 8'hf4 : _GEN_1465; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1467 = 8'hbb == inBytes_5 ? 8'hea : _GEN_1466; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1468 = 8'hbc == inBytes_5 ? 8'h65 : _GEN_1467; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1469 = 8'hbd == inBytes_5 ? 8'h7a : _GEN_1468; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1470 = 8'hbe == inBytes_5 ? 8'hae : _GEN_1469; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1471 = 8'hbf == inBytes_5 ? 8'h8 : _GEN_1470; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1472 = 8'hc0 == inBytes_5 ? 8'hba : _GEN_1471; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1473 = 8'hc1 == inBytes_5 ? 8'h78 : _GEN_1472; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1474 = 8'hc2 == inBytes_5 ? 8'h25 : _GEN_1473; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1475 = 8'hc3 == inBytes_5 ? 8'h2e : _GEN_1474; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1476 = 8'hc4 == inBytes_5 ? 8'h1c : _GEN_1475; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1477 = 8'hc5 == inBytes_5 ? 8'ha6 : _GEN_1476; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1478 = 8'hc6 == inBytes_5 ? 8'hb4 : _GEN_1477; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1479 = 8'hc7 == inBytes_5 ? 8'hc6 : _GEN_1478; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1480 = 8'hc8 == inBytes_5 ? 8'he8 : _GEN_1479; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1481 = 8'hc9 == inBytes_5 ? 8'hdd : _GEN_1480; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1482 = 8'hca == inBytes_5 ? 8'h74 : _GEN_1481; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1483 = 8'hcb == inBytes_5 ? 8'h1f : _GEN_1482; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1484 = 8'hcc == inBytes_5 ? 8'h4b : _GEN_1483; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1485 = 8'hcd == inBytes_5 ? 8'hbd : _GEN_1484; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1486 = 8'hce == inBytes_5 ? 8'h8b : _GEN_1485; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1487 = 8'hcf == inBytes_5 ? 8'h8a : _GEN_1486; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1488 = 8'hd0 == inBytes_5 ? 8'h70 : _GEN_1487; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1489 = 8'hd1 == inBytes_5 ? 8'h3e : _GEN_1488; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1490 = 8'hd2 == inBytes_5 ? 8'hb5 : _GEN_1489; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1491 = 8'hd3 == inBytes_5 ? 8'h66 : _GEN_1490; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1492 = 8'hd4 == inBytes_5 ? 8'h48 : _GEN_1491; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1493 = 8'hd5 == inBytes_5 ? 8'h3 : _GEN_1492; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1494 = 8'hd6 == inBytes_5 ? 8'hf6 : _GEN_1493; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1495 = 8'hd7 == inBytes_5 ? 8'he : _GEN_1494; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1496 = 8'hd8 == inBytes_5 ? 8'h61 : _GEN_1495; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1497 = 8'hd9 == inBytes_5 ? 8'h35 : _GEN_1496; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1498 = 8'hda == inBytes_5 ? 8'h57 : _GEN_1497; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1499 = 8'hdb == inBytes_5 ? 8'hb9 : _GEN_1498; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1500 = 8'hdc == inBytes_5 ? 8'h86 : _GEN_1499; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1501 = 8'hdd == inBytes_5 ? 8'hc1 : _GEN_1500; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1502 = 8'hde == inBytes_5 ? 8'h1d : _GEN_1501; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1503 = 8'hdf == inBytes_5 ? 8'h9e : _GEN_1502; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1504 = 8'he0 == inBytes_5 ? 8'he1 : _GEN_1503; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1505 = 8'he1 == inBytes_5 ? 8'hf8 : _GEN_1504; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1506 = 8'he2 == inBytes_5 ? 8'h98 : _GEN_1505; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1507 = 8'he3 == inBytes_5 ? 8'h11 : _GEN_1506; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1508 = 8'he4 == inBytes_5 ? 8'h69 : _GEN_1507; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1509 = 8'he5 == inBytes_5 ? 8'hd9 : _GEN_1508; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1510 = 8'he6 == inBytes_5 ? 8'h8e : _GEN_1509; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1511 = 8'he7 == inBytes_5 ? 8'h94 : _GEN_1510; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1512 = 8'he8 == inBytes_5 ? 8'h9b : _GEN_1511; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1513 = 8'he9 == inBytes_5 ? 8'h1e : _GEN_1512; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1514 = 8'hea == inBytes_5 ? 8'h87 : _GEN_1513; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1515 = 8'heb == inBytes_5 ? 8'he9 : _GEN_1514; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1516 = 8'hec == inBytes_5 ? 8'hce : _GEN_1515; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1517 = 8'hed == inBytes_5 ? 8'h55 : _GEN_1516; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1518 = 8'hee == inBytes_5 ? 8'h28 : _GEN_1517; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1519 = 8'hef == inBytes_5 ? 8'hdf : _GEN_1518; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1520 = 8'hf0 == inBytes_5 ? 8'h8c : _GEN_1519; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1521 = 8'hf1 == inBytes_5 ? 8'ha1 : _GEN_1520; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1522 = 8'hf2 == inBytes_5 ? 8'h89 : _GEN_1521; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1523 = 8'hf3 == inBytes_5 ? 8'hd : _GEN_1522; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1524 = 8'hf4 == inBytes_5 ? 8'hbf : _GEN_1523; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1525 = 8'hf5 == inBytes_5 ? 8'he6 : _GEN_1524; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1526 = 8'hf6 == inBytes_5 ? 8'h42 : _GEN_1525; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1527 = 8'hf7 == inBytes_5 ? 8'h68 : _GEN_1526; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1528 = 8'hf8 == inBytes_5 ? 8'h41 : _GEN_1527; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1529 = 8'hf9 == inBytes_5 ? 8'h99 : _GEN_1528; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1530 = 8'hfa == inBytes_5 ? 8'h2d : _GEN_1529; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1531 = 8'hfb == inBytes_5 ? 8'hf : _GEN_1530; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1532 = 8'hfc == inBytes_5 ? 8'hb0 : _GEN_1531; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1533 = 8'hfd == inBytes_5 ? 8'h54 : _GEN_1532; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1534 = 8'hfe == inBytes_5 ? 8'hbb : _GEN_1533; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] outBytes_5 = 8'hff == inBytes_5 ? 8'h16 : _GEN_1534; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1537 = 8'h1 == inBytes_6 ? 8'h7c : 8'h63; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1538 = 8'h2 == inBytes_6 ? 8'h77 : _GEN_1537; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1539 = 8'h3 == inBytes_6 ? 8'h7b : _GEN_1538; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1540 = 8'h4 == inBytes_6 ? 8'hf2 : _GEN_1539; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1541 = 8'h5 == inBytes_6 ? 8'h6b : _GEN_1540; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1542 = 8'h6 == inBytes_6 ? 8'h6f : _GEN_1541; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1543 = 8'h7 == inBytes_6 ? 8'hc5 : _GEN_1542; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1544 = 8'h8 == inBytes_6 ? 8'h30 : _GEN_1543; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1545 = 8'h9 == inBytes_6 ? 8'h1 : _GEN_1544; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1546 = 8'ha == inBytes_6 ? 8'h67 : _GEN_1545; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1547 = 8'hb == inBytes_6 ? 8'h2b : _GEN_1546; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1548 = 8'hc == inBytes_6 ? 8'hfe : _GEN_1547; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1549 = 8'hd == inBytes_6 ? 8'hd7 : _GEN_1548; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1550 = 8'he == inBytes_6 ? 8'hab : _GEN_1549; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1551 = 8'hf == inBytes_6 ? 8'h76 : _GEN_1550; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1552 = 8'h10 == inBytes_6 ? 8'hca : _GEN_1551; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1553 = 8'h11 == inBytes_6 ? 8'h82 : _GEN_1552; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1554 = 8'h12 == inBytes_6 ? 8'hc9 : _GEN_1553; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1555 = 8'h13 == inBytes_6 ? 8'h7d : _GEN_1554; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1556 = 8'h14 == inBytes_6 ? 8'hfa : _GEN_1555; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1557 = 8'h15 == inBytes_6 ? 8'h59 : _GEN_1556; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1558 = 8'h16 == inBytes_6 ? 8'h47 : _GEN_1557; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1559 = 8'h17 == inBytes_6 ? 8'hf0 : _GEN_1558; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1560 = 8'h18 == inBytes_6 ? 8'had : _GEN_1559; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1561 = 8'h19 == inBytes_6 ? 8'hd4 : _GEN_1560; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1562 = 8'h1a == inBytes_6 ? 8'ha2 : _GEN_1561; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1563 = 8'h1b == inBytes_6 ? 8'haf : _GEN_1562; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1564 = 8'h1c == inBytes_6 ? 8'h9c : _GEN_1563; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1565 = 8'h1d == inBytes_6 ? 8'ha4 : _GEN_1564; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1566 = 8'h1e == inBytes_6 ? 8'h72 : _GEN_1565; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1567 = 8'h1f == inBytes_6 ? 8'hc0 : _GEN_1566; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1568 = 8'h20 == inBytes_6 ? 8'hb7 : _GEN_1567; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1569 = 8'h21 == inBytes_6 ? 8'hfd : _GEN_1568; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1570 = 8'h22 == inBytes_6 ? 8'h93 : _GEN_1569; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1571 = 8'h23 == inBytes_6 ? 8'h26 : _GEN_1570; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1572 = 8'h24 == inBytes_6 ? 8'h36 : _GEN_1571; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1573 = 8'h25 == inBytes_6 ? 8'h3f : _GEN_1572; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1574 = 8'h26 == inBytes_6 ? 8'hf7 : _GEN_1573; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1575 = 8'h27 == inBytes_6 ? 8'hcc : _GEN_1574; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1576 = 8'h28 == inBytes_6 ? 8'h34 : _GEN_1575; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1577 = 8'h29 == inBytes_6 ? 8'ha5 : _GEN_1576; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1578 = 8'h2a == inBytes_6 ? 8'he5 : _GEN_1577; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1579 = 8'h2b == inBytes_6 ? 8'hf1 : _GEN_1578; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1580 = 8'h2c == inBytes_6 ? 8'h71 : _GEN_1579; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1581 = 8'h2d == inBytes_6 ? 8'hd8 : _GEN_1580; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1582 = 8'h2e == inBytes_6 ? 8'h31 : _GEN_1581; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1583 = 8'h2f == inBytes_6 ? 8'h15 : _GEN_1582; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1584 = 8'h30 == inBytes_6 ? 8'h4 : _GEN_1583; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1585 = 8'h31 == inBytes_6 ? 8'hc7 : _GEN_1584; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1586 = 8'h32 == inBytes_6 ? 8'h23 : _GEN_1585; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1587 = 8'h33 == inBytes_6 ? 8'hc3 : _GEN_1586; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1588 = 8'h34 == inBytes_6 ? 8'h18 : _GEN_1587; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1589 = 8'h35 == inBytes_6 ? 8'h96 : _GEN_1588; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1590 = 8'h36 == inBytes_6 ? 8'h5 : _GEN_1589; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1591 = 8'h37 == inBytes_6 ? 8'h9a : _GEN_1590; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1592 = 8'h38 == inBytes_6 ? 8'h7 : _GEN_1591; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1593 = 8'h39 == inBytes_6 ? 8'h12 : _GEN_1592; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1594 = 8'h3a == inBytes_6 ? 8'h80 : _GEN_1593; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1595 = 8'h3b == inBytes_6 ? 8'he2 : _GEN_1594; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1596 = 8'h3c == inBytes_6 ? 8'heb : _GEN_1595; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1597 = 8'h3d == inBytes_6 ? 8'h27 : _GEN_1596; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1598 = 8'h3e == inBytes_6 ? 8'hb2 : _GEN_1597; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1599 = 8'h3f == inBytes_6 ? 8'h75 : _GEN_1598; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1600 = 8'h40 == inBytes_6 ? 8'h9 : _GEN_1599; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1601 = 8'h41 == inBytes_6 ? 8'h83 : _GEN_1600; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1602 = 8'h42 == inBytes_6 ? 8'h2c : _GEN_1601; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1603 = 8'h43 == inBytes_6 ? 8'h1a : _GEN_1602; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1604 = 8'h44 == inBytes_6 ? 8'h1b : _GEN_1603; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1605 = 8'h45 == inBytes_6 ? 8'h6e : _GEN_1604; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1606 = 8'h46 == inBytes_6 ? 8'h5a : _GEN_1605; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1607 = 8'h47 == inBytes_6 ? 8'ha0 : _GEN_1606; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1608 = 8'h48 == inBytes_6 ? 8'h52 : _GEN_1607; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1609 = 8'h49 == inBytes_6 ? 8'h3b : _GEN_1608; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1610 = 8'h4a == inBytes_6 ? 8'hd6 : _GEN_1609; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1611 = 8'h4b == inBytes_6 ? 8'hb3 : _GEN_1610; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1612 = 8'h4c == inBytes_6 ? 8'h29 : _GEN_1611; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1613 = 8'h4d == inBytes_6 ? 8'he3 : _GEN_1612; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1614 = 8'h4e == inBytes_6 ? 8'h2f : _GEN_1613; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1615 = 8'h4f == inBytes_6 ? 8'h84 : _GEN_1614; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1616 = 8'h50 == inBytes_6 ? 8'h53 : _GEN_1615; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1617 = 8'h51 == inBytes_6 ? 8'hd1 : _GEN_1616; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1618 = 8'h52 == inBytes_6 ? 8'h0 : _GEN_1617; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1619 = 8'h53 == inBytes_6 ? 8'hed : _GEN_1618; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1620 = 8'h54 == inBytes_6 ? 8'h20 : _GEN_1619; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1621 = 8'h55 == inBytes_6 ? 8'hfc : _GEN_1620; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1622 = 8'h56 == inBytes_6 ? 8'hb1 : _GEN_1621; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1623 = 8'h57 == inBytes_6 ? 8'h5b : _GEN_1622; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1624 = 8'h58 == inBytes_6 ? 8'h6a : _GEN_1623; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1625 = 8'h59 == inBytes_6 ? 8'hcb : _GEN_1624; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1626 = 8'h5a == inBytes_6 ? 8'hbe : _GEN_1625; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1627 = 8'h5b == inBytes_6 ? 8'h39 : _GEN_1626; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1628 = 8'h5c == inBytes_6 ? 8'h4a : _GEN_1627; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1629 = 8'h5d == inBytes_6 ? 8'h4c : _GEN_1628; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1630 = 8'h5e == inBytes_6 ? 8'h58 : _GEN_1629; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1631 = 8'h5f == inBytes_6 ? 8'hcf : _GEN_1630; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1632 = 8'h60 == inBytes_6 ? 8'hd0 : _GEN_1631; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1633 = 8'h61 == inBytes_6 ? 8'hef : _GEN_1632; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1634 = 8'h62 == inBytes_6 ? 8'haa : _GEN_1633; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1635 = 8'h63 == inBytes_6 ? 8'hfb : _GEN_1634; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1636 = 8'h64 == inBytes_6 ? 8'h43 : _GEN_1635; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1637 = 8'h65 == inBytes_6 ? 8'h4d : _GEN_1636; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1638 = 8'h66 == inBytes_6 ? 8'h33 : _GEN_1637; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1639 = 8'h67 == inBytes_6 ? 8'h85 : _GEN_1638; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1640 = 8'h68 == inBytes_6 ? 8'h45 : _GEN_1639; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1641 = 8'h69 == inBytes_6 ? 8'hf9 : _GEN_1640; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1642 = 8'h6a == inBytes_6 ? 8'h2 : _GEN_1641; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1643 = 8'h6b == inBytes_6 ? 8'h7f : _GEN_1642; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1644 = 8'h6c == inBytes_6 ? 8'h50 : _GEN_1643; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1645 = 8'h6d == inBytes_6 ? 8'h3c : _GEN_1644; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1646 = 8'h6e == inBytes_6 ? 8'h9f : _GEN_1645; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1647 = 8'h6f == inBytes_6 ? 8'ha8 : _GEN_1646; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1648 = 8'h70 == inBytes_6 ? 8'h51 : _GEN_1647; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1649 = 8'h71 == inBytes_6 ? 8'ha3 : _GEN_1648; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1650 = 8'h72 == inBytes_6 ? 8'h40 : _GEN_1649; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1651 = 8'h73 == inBytes_6 ? 8'h8f : _GEN_1650; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1652 = 8'h74 == inBytes_6 ? 8'h92 : _GEN_1651; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1653 = 8'h75 == inBytes_6 ? 8'h9d : _GEN_1652; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1654 = 8'h76 == inBytes_6 ? 8'h38 : _GEN_1653; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1655 = 8'h77 == inBytes_6 ? 8'hf5 : _GEN_1654; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1656 = 8'h78 == inBytes_6 ? 8'hbc : _GEN_1655; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1657 = 8'h79 == inBytes_6 ? 8'hb6 : _GEN_1656; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1658 = 8'h7a == inBytes_6 ? 8'hda : _GEN_1657; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1659 = 8'h7b == inBytes_6 ? 8'h21 : _GEN_1658; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1660 = 8'h7c == inBytes_6 ? 8'h10 : _GEN_1659; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1661 = 8'h7d == inBytes_6 ? 8'hff : _GEN_1660; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1662 = 8'h7e == inBytes_6 ? 8'hf3 : _GEN_1661; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1663 = 8'h7f == inBytes_6 ? 8'hd2 : _GEN_1662; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1664 = 8'h80 == inBytes_6 ? 8'hcd : _GEN_1663; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1665 = 8'h81 == inBytes_6 ? 8'hc : _GEN_1664; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1666 = 8'h82 == inBytes_6 ? 8'h13 : _GEN_1665; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1667 = 8'h83 == inBytes_6 ? 8'hec : _GEN_1666; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1668 = 8'h84 == inBytes_6 ? 8'h5f : _GEN_1667; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1669 = 8'h85 == inBytes_6 ? 8'h97 : _GEN_1668; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1670 = 8'h86 == inBytes_6 ? 8'h44 : _GEN_1669; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1671 = 8'h87 == inBytes_6 ? 8'h17 : _GEN_1670; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1672 = 8'h88 == inBytes_6 ? 8'hc4 : _GEN_1671; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1673 = 8'h89 == inBytes_6 ? 8'ha7 : _GEN_1672; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1674 = 8'h8a == inBytes_6 ? 8'h7e : _GEN_1673; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1675 = 8'h8b == inBytes_6 ? 8'h3d : _GEN_1674; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1676 = 8'h8c == inBytes_6 ? 8'h64 : _GEN_1675; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1677 = 8'h8d == inBytes_6 ? 8'h5d : _GEN_1676; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1678 = 8'h8e == inBytes_6 ? 8'h19 : _GEN_1677; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1679 = 8'h8f == inBytes_6 ? 8'h73 : _GEN_1678; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1680 = 8'h90 == inBytes_6 ? 8'h60 : _GEN_1679; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1681 = 8'h91 == inBytes_6 ? 8'h81 : _GEN_1680; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1682 = 8'h92 == inBytes_6 ? 8'h4f : _GEN_1681; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1683 = 8'h93 == inBytes_6 ? 8'hdc : _GEN_1682; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1684 = 8'h94 == inBytes_6 ? 8'h22 : _GEN_1683; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1685 = 8'h95 == inBytes_6 ? 8'h2a : _GEN_1684; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1686 = 8'h96 == inBytes_6 ? 8'h90 : _GEN_1685; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1687 = 8'h97 == inBytes_6 ? 8'h88 : _GEN_1686; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1688 = 8'h98 == inBytes_6 ? 8'h46 : _GEN_1687; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1689 = 8'h99 == inBytes_6 ? 8'hee : _GEN_1688; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1690 = 8'h9a == inBytes_6 ? 8'hb8 : _GEN_1689; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1691 = 8'h9b == inBytes_6 ? 8'h14 : _GEN_1690; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1692 = 8'h9c == inBytes_6 ? 8'hde : _GEN_1691; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1693 = 8'h9d == inBytes_6 ? 8'h5e : _GEN_1692; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1694 = 8'h9e == inBytes_6 ? 8'hb : _GEN_1693; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1695 = 8'h9f == inBytes_6 ? 8'hdb : _GEN_1694; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1696 = 8'ha0 == inBytes_6 ? 8'he0 : _GEN_1695; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1697 = 8'ha1 == inBytes_6 ? 8'h32 : _GEN_1696; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1698 = 8'ha2 == inBytes_6 ? 8'h3a : _GEN_1697; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1699 = 8'ha3 == inBytes_6 ? 8'ha : _GEN_1698; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1700 = 8'ha4 == inBytes_6 ? 8'h49 : _GEN_1699; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1701 = 8'ha5 == inBytes_6 ? 8'h6 : _GEN_1700; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1702 = 8'ha6 == inBytes_6 ? 8'h24 : _GEN_1701; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1703 = 8'ha7 == inBytes_6 ? 8'h5c : _GEN_1702; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1704 = 8'ha8 == inBytes_6 ? 8'hc2 : _GEN_1703; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1705 = 8'ha9 == inBytes_6 ? 8'hd3 : _GEN_1704; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1706 = 8'haa == inBytes_6 ? 8'hac : _GEN_1705; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1707 = 8'hab == inBytes_6 ? 8'h62 : _GEN_1706; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1708 = 8'hac == inBytes_6 ? 8'h91 : _GEN_1707; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1709 = 8'had == inBytes_6 ? 8'h95 : _GEN_1708; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1710 = 8'hae == inBytes_6 ? 8'he4 : _GEN_1709; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1711 = 8'haf == inBytes_6 ? 8'h79 : _GEN_1710; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1712 = 8'hb0 == inBytes_6 ? 8'he7 : _GEN_1711; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1713 = 8'hb1 == inBytes_6 ? 8'hc8 : _GEN_1712; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1714 = 8'hb2 == inBytes_6 ? 8'h37 : _GEN_1713; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1715 = 8'hb3 == inBytes_6 ? 8'h6d : _GEN_1714; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1716 = 8'hb4 == inBytes_6 ? 8'h8d : _GEN_1715; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1717 = 8'hb5 == inBytes_6 ? 8'hd5 : _GEN_1716; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1718 = 8'hb6 == inBytes_6 ? 8'h4e : _GEN_1717; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1719 = 8'hb7 == inBytes_6 ? 8'ha9 : _GEN_1718; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1720 = 8'hb8 == inBytes_6 ? 8'h6c : _GEN_1719; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1721 = 8'hb9 == inBytes_6 ? 8'h56 : _GEN_1720; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1722 = 8'hba == inBytes_6 ? 8'hf4 : _GEN_1721; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1723 = 8'hbb == inBytes_6 ? 8'hea : _GEN_1722; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1724 = 8'hbc == inBytes_6 ? 8'h65 : _GEN_1723; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1725 = 8'hbd == inBytes_6 ? 8'h7a : _GEN_1724; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1726 = 8'hbe == inBytes_6 ? 8'hae : _GEN_1725; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1727 = 8'hbf == inBytes_6 ? 8'h8 : _GEN_1726; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1728 = 8'hc0 == inBytes_6 ? 8'hba : _GEN_1727; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1729 = 8'hc1 == inBytes_6 ? 8'h78 : _GEN_1728; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1730 = 8'hc2 == inBytes_6 ? 8'h25 : _GEN_1729; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1731 = 8'hc3 == inBytes_6 ? 8'h2e : _GEN_1730; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1732 = 8'hc4 == inBytes_6 ? 8'h1c : _GEN_1731; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1733 = 8'hc5 == inBytes_6 ? 8'ha6 : _GEN_1732; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1734 = 8'hc6 == inBytes_6 ? 8'hb4 : _GEN_1733; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1735 = 8'hc7 == inBytes_6 ? 8'hc6 : _GEN_1734; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1736 = 8'hc8 == inBytes_6 ? 8'he8 : _GEN_1735; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1737 = 8'hc9 == inBytes_6 ? 8'hdd : _GEN_1736; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1738 = 8'hca == inBytes_6 ? 8'h74 : _GEN_1737; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1739 = 8'hcb == inBytes_6 ? 8'h1f : _GEN_1738; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1740 = 8'hcc == inBytes_6 ? 8'h4b : _GEN_1739; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1741 = 8'hcd == inBytes_6 ? 8'hbd : _GEN_1740; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1742 = 8'hce == inBytes_6 ? 8'h8b : _GEN_1741; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1743 = 8'hcf == inBytes_6 ? 8'h8a : _GEN_1742; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1744 = 8'hd0 == inBytes_6 ? 8'h70 : _GEN_1743; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1745 = 8'hd1 == inBytes_6 ? 8'h3e : _GEN_1744; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1746 = 8'hd2 == inBytes_6 ? 8'hb5 : _GEN_1745; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1747 = 8'hd3 == inBytes_6 ? 8'h66 : _GEN_1746; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1748 = 8'hd4 == inBytes_6 ? 8'h48 : _GEN_1747; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1749 = 8'hd5 == inBytes_6 ? 8'h3 : _GEN_1748; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1750 = 8'hd6 == inBytes_6 ? 8'hf6 : _GEN_1749; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1751 = 8'hd7 == inBytes_6 ? 8'he : _GEN_1750; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1752 = 8'hd8 == inBytes_6 ? 8'h61 : _GEN_1751; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1753 = 8'hd9 == inBytes_6 ? 8'h35 : _GEN_1752; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1754 = 8'hda == inBytes_6 ? 8'h57 : _GEN_1753; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1755 = 8'hdb == inBytes_6 ? 8'hb9 : _GEN_1754; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1756 = 8'hdc == inBytes_6 ? 8'h86 : _GEN_1755; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1757 = 8'hdd == inBytes_6 ? 8'hc1 : _GEN_1756; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1758 = 8'hde == inBytes_6 ? 8'h1d : _GEN_1757; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1759 = 8'hdf == inBytes_6 ? 8'h9e : _GEN_1758; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1760 = 8'he0 == inBytes_6 ? 8'he1 : _GEN_1759; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1761 = 8'he1 == inBytes_6 ? 8'hf8 : _GEN_1760; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1762 = 8'he2 == inBytes_6 ? 8'h98 : _GEN_1761; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1763 = 8'he3 == inBytes_6 ? 8'h11 : _GEN_1762; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1764 = 8'he4 == inBytes_6 ? 8'h69 : _GEN_1763; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1765 = 8'he5 == inBytes_6 ? 8'hd9 : _GEN_1764; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1766 = 8'he6 == inBytes_6 ? 8'h8e : _GEN_1765; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1767 = 8'he7 == inBytes_6 ? 8'h94 : _GEN_1766; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1768 = 8'he8 == inBytes_6 ? 8'h9b : _GEN_1767; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1769 = 8'he9 == inBytes_6 ? 8'h1e : _GEN_1768; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1770 = 8'hea == inBytes_6 ? 8'h87 : _GEN_1769; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1771 = 8'heb == inBytes_6 ? 8'he9 : _GEN_1770; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1772 = 8'hec == inBytes_6 ? 8'hce : _GEN_1771; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1773 = 8'hed == inBytes_6 ? 8'h55 : _GEN_1772; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1774 = 8'hee == inBytes_6 ? 8'h28 : _GEN_1773; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1775 = 8'hef == inBytes_6 ? 8'hdf : _GEN_1774; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1776 = 8'hf0 == inBytes_6 ? 8'h8c : _GEN_1775; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1777 = 8'hf1 == inBytes_6 ? 8'ha1 : _GEN_1776; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1778 = 8'hf2 == inBytes_6 ? 8'h89 : _GEN_1777; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1779 = 8'hf3 == inBytes_6 ? 8'hd : _GEN_1778; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1780 = 8'hf4 == inBytes_6 ? 8'hbf : _GEN_1779; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1781 = 8'hf5 == inBytes_6 ? 8'he6 : _GEN_1780; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1782 = 8'hf6 == inBytes_6 ? 8'h42 : _GEN_1781; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1783 = 8'hf7 == inBytes_6 ? 8'h68 : _GEN_1782; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1784 = 8'hf8 == inBytes_6 ? 8'h41 : _GEN_1783; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1785 = 8'hf9 == inBytes_6 ? 8'h99 : _GEN_1784; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1786 = 8'hfa == inBytes_6 ? 8'h2d : _GEN_1785; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1787 = 8'hfb == inBytes_6 ? 8'hf : _GEN_1786; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1788 = 8'hfc == inBytes_6 ? 8'hb0 : _GEN_1787; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1789 = 8'hfd == inBytes_6 ? 8'h54 : _GEN_1788; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1790 = 8'hfe == inBytes_6 ? 8'hbb : _GEN_1789; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] outBytes_6 = 8'hff == inBytes_6 ? 8'h16 : _GEN_1790; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1793 = 8'h1 == inBytes_7 ? 8'h7c : 8'h63; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1794 = 8'h2 == inBytes_7 ? 8'h77 : _GEN_1793; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1795 = 8'h3 == inBytes_7 ? 8'h7b : _GEN_1794; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1796 = 8'h4 == inBytes_7 ? 8'hf2 : _GEN_1795; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1797 = 8'h5 == inBytes_7 ? 8'h6b : _GEN_1796; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1798 = 8'h6 == inBytes_7 ? 8'h6f : _GEN_1797; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1799 = 8'h7 == inBytes_7 ? 8'hc5 : _GEN_1798; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1800 = 8'h8 == inBytes_7 ? 8'h30 : _GEN_1799; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1801 = 8'h9 == inBytes_7 ? 8'h1 : _GEN_1800; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1802 = 8'ha == inBytes_7 ? 8'h67 : _GEN_1801; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1803 = 8'hb == inBytes_7 ? 8'h2b : _GEN_1802; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1804 = 8'hc == inBytes_7 ? 8'hfe : _GEN_1803; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1805 = 8'hd == inBytes_7 ? 8'hd7 : _GEN_1804; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1806 = 8'he == inBytes_7 ? 8'hab : _GEN_1805; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1807 = 8'hf == inBytes_7 ? 8'h76 : _GEN_1806; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1808 = 8'h10 == inBytes_7 ? 8'hca : _GEN_1807; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1809 = 8'h11 == inBytes_7 ? 8'h82 : _GEN_1808; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1810 = 8'h12 == inBytes_7 ? 8'hc9 : _GEN_1809; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1811 = 8'h13 == inBytes_7 ? 8'h7d : _GEN_1810; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1812 = 8'h14 == inBytes_7 ? 8'hfa : _GEN_1811; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1813 = 8'h15 == inBytes_7 ? 8'h59 : _GEN_1812; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1814 = 8'h16 == inBytes_7 ? 8'h47 : _GEN_1813; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1815 = 8'h17 == inBytes_7 ? 8'hf0 : _GEN_1814; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1816 = 8'h18 == inBytes_7 ? 8'had : _GEN_1815; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1817 = 8'h19 == inBytes_7 ? 8'hd4 : _GEN_1816; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1818 = 8'h1a == inBytes_7 ? 8'ha2 : _GEN_1817; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1819 = 8'h1b == inBytes_7 ? 8'haf : _GEN_1818; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1820 = 8'h1c == inBytes_7 ? 8'h9c : _GEN_1819; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1821 = 8'h1d == inBytes_7 ? 8'ha4 : _GEN_1820; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1822 = 8'h1e == inBytes_7 ? 8'h72 : _GEN_1821; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1823 = 8'h1f == inBytes_7 ? 8'hc0 : _GEN_1822; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1824 = 8'h20 == inBytes_7 ? 8'hb7 : _GEN_1823; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1825 = 8'h21 == inBytes_7 ? 8'hfd : _GEN_1824; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1826 = 8'h22 == inBytes_7 ? 8'h93 : _GEN_1825; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1827 = 8'h23 == inBytes_7 ? 8'h26 : _GEN_1826; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1828 = 8'h24 == inBytes_7 ? 8'h36 : _GEN_1827; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1829 = 8'h25 == inBytes_7 ? 8'h3f : _GEN_1828; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1830 = 8'h26 == inBytes_7 ? 8'hf7 : _GEN_1829; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1831 = 8'h27 == inBytes_7 ? 8'hcc : _GEN_1830; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1832 = 8'h28 == inBytes_7 ? 8'h34 : _GEN_1831; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1833 = 8'h29 == inBytes_7 ? 8'ha5 : _GEN_1832; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1834 = 8'h2a == inBytes_7 ? 8'he5 : _GEN_1833; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1835 = 8'h2b == inBytes_7 ? 8'hf1 : _GEN_1834; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1836 = 8'h2c == inBytes_7 ? 8'h71 : _GEN_1835; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1837 = 8'h2d == inBytes_7 ? 8'hd8 : _GEN_1836; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1838 = 8'h2e == inBytes_7 ? 8'h31 : _GEN_1837; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1839 = 8'h2f == inBytes_7 ? 8'h15 : _GEN_1838; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1840 = 8'h30 == inBytes_7 ? 8'h4 : _GEN_1839; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1841 = 8'h31 == inBytes_7 ? 8'hc7 : _GEN_1840; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1842 = 8'h32 == inBytes_7 ? 8'h23 : _GEN_1841; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1843 = 8'h33 == inBytes_7 ? 8'hc3 : _GEN_1842; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1844 = 8'h34 == inBytes_7 ? 8'h18 : _GEN_1843; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1845 = 8'h35 == inBytes_7 ? 8'h96 : _GEN_1844; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1846 = 8'h36 == inBytes_7 ? 8'h5 : _GEN_1845; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1847 = 8'h37 == inBytes_7 ? 8'h9a : _GEN_1846; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1848 = 8'h38 == inBytes_7 ? 8'h7 : _GEN_1847; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1849 = 8'h39 == inBytes_7 ? 8'h12 : _GEN_1848; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1850 = 8'h3a == inBytes_7 ? 8'h80 : _GEN_1849; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1851 = 8'h3b == inBytes_7 ? 8'he2 : _GEN_1850; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1852 = 8'h3c == inBytes_7 ? 8'heb : _GEN_1851; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1853 = 8'h3d == inBytes_7 ? 8'h27 : _GEN_1852; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1854 = 8'h3e == inBytes_7 ? 8'hb2 : _GEN_1853; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1855 = 8'h3f == inBytes_7 ? 8'h75 : _GEN_1854; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1856 = 8'h40 == inBytes_7 ? 8'h9 : _GEN_1855; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1857 = 8'h41 == inBytes_7 ? 8'h83 : _GEN_1856; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1858 = 8'h42 == inBytes_7 ? 8'h2c : _GEN_1857; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1859 = 8'h43 == inBytes_7 ? 8'h1a : _GEN_1858; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1860 = 8'h44 == inBytes_7 ? 8'h1b : _GEN_1859; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1861 = 8'h45 == inBytes_7 ? 8'h6e : _GEN_1860; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1862 = 8'h46 == inBytes_7 ? 8'h5a : _GEN_1861; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1863 = 8'h47 == inBytes_7 ? 8'ha0 : _GEN_1862; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1864 = 8'h48 == inBytes_7 ? 8'h52 : _GEN_1863; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1865 = 8'h49 == inBytes_7 ? 8'h3b : _GEN_1864; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1866 = 8'h4a == inBytes_7 ? 8'hd6 : _GEN_1865; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1867 = 8'h4b == inBytes_7 ? 8'hb3 : _GEN_1866; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1868 = 8'h4c == inBytes_7 ? 8'h29 : _GEN_1867; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1869 = 8'h4d == inBytes_7 ? 8'he3 : _GEN_1868; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1870 = 8'h4e == inBytes_7 ? 8'h2f : _GEN_1869; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1871 = 8'h4f == inBytes_7 ? 8'h84 : _GEN_1870; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1872 = 8'h50 == inBytes_7 ? 8'h53 : _GEN_1871; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1873 = 8'h51 == inBytes_7 ? 8'hd1 : _GEN_1872; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1874 = 8'h52 == inBytes_7 ? 8'h0 : _GEN_1873; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1875 = 8'h53 == inBytes_7 ? 8'hed : _GEN_1874; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1876 = 8'h54 == inBytes_7 ? 8'h20 : _GEN_1875; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1877 = 8'h55 == inBytes_7 ? 8'hfc : _GEN_1876; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1878 = 8'h56 == inBytes_7 ? 8'hb1 : _GEN_1877; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1879 = 8'h57 == inBytes_7 ? 8'h5b : _GEN_1878; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1880 = 8'h58 == inBytes_7 ? 8'h6a : _GEN_1879; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1881 = 8'h59 == inBytes_7 ? 8'hcb : _GEN_1880; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1882 = 8'h5a == inBytes_7 ? 8'hbe : _GEN_1881; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1883 = 8'h5b == inBytes_7 ? 8'h39 : _GEN_1882; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1884 = 8'h5c == inBytes_7 ? 8'h4a : _GEN_1883; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1885 = 8'h5d == inBytes_7 ? 8'h4c : _GEN_1884; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1886 = 8'h5e == inBytes_7 ? 8'h58 : _GEN_1885; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1887 = 8'h5f == inBytes_7 ? 8'hcf : _GEN_1886; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1888 = 8'h60 == inBytes_7 ? 8'hd0 : _GEN_1887; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1889 = 8'h61 == inBytes_7 ? 8'hef : _GEN_1888; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1890 = 8'h62 == inBytes_7 ? 8'haa : _GEN_1889; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1891 = 8'h63 == inBytes_7 ? 8'hfb : _GEN_1890; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1892 = 8'h64 == inBytes_7 ? 8'h43 : _GEN_1891; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1893 = 8'h65 == inBytes_7 ? 8'h4d : _GEN_1892; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1894 = 8'h66 == inBytes_7 ? 8'h33 : _GEN_1893; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1895 = 8'h67 == inBytes_7 ? 8'h85 : _GEN_1894; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1896 = 8'h68 == inBytes_7 ? 8'h45 : _GEN_1895; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1897 = 8'h69 == inBytes_7 ? 8'hf9 : _GEN_1896; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1898 = 8'h6a == inBytes_7 ? 8'h2 : _GEN_1897; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1899 = 8'h6b == inBytes_7 ? 8'h7f : _GEN_1898; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1900 = 8'h6c == inBytes_7 ? 8'h50 : _GEN_1899; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1901 = 8'h6d == inBytes_7 ? 8'h3c : _GEN_1900; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1902 = 8'h6e == inBytes_7 ? 8'h9f : _GEN_1901; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1903 = 8'h6f == inBytes_7 ? 8'ha8 : _GEN_1902; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1904 = 8'h70 == inBytes_7 ? 8'h51 : _GEN_1903; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1905 = 8'h71 == inBytes_7 ? 8'ha3 : _GEN_1904; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1906 = 8'h72 == inBytes_7 ? 8'h40 : _GEN_1905; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1907 = 8'h73 == inBytes_7 ? 8'h8f : _GEN_1906; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1908 = 8'h74 == inBytes_7 ? 8'h92 : _GEN_1907; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1909 = 8'h75 == inBytes_7 ? 8'h9d : _GEN_1908; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1910 = 8'h76 == inBytes_7 ? 8'h38 : _GEN_1909; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1911 = 8'h77 == inBytes_7 ? 8'hf5 : _GEN_1910; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1912 = 8'h78 == inBytes_7 ? 8'hbc : _GEN_1911; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1913 = 8'h79 == inBytes_7 ? 8'hb6 : _GEN_1912; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1914 = 8'h7a == inBytes_7 ? 8'hda : _GEN_1913; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1915 = 8'h7b == inBytes_7 ? 8'h21 : _GEN_1914; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1916 = 8'h7c == inBytes_7 ? 8'h10 : _GEN_1915; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1917 = 8'h7d == inBytes_7 ? 8'hff : _GEN_1916; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1918 = 8'h7e == inBytes_7 ? 8'hf3 : _GEN_1917; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1919 = 8'h7f == inBytes_7 ? 8'hd2 : _GEN_1918; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1920 = 8'h80 == inBytes_7 ? 8'hcd : _GEN_1919; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1921 = 8'h81 == inBytes_7 ? 8'hc : _GEN_1920; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1922 = 8'h82 == inBytes_7 ? 8'h13 : _GEN_1921; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1923 = 8'h83 == inBytes_7 ? 8'hec : _GEN_1922; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1924 = 8'h84 == inBytes_7 ? 8'h5f : _GEN_1923; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1925 = 8'h85 == inBytes_7 ? 8'h97 : _GEN_1924; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1926 = 8'h86 == inBytes_7 ? 8'h44 : _GEN_1925; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1927 = 8'h87 == inBytes_7 ? 8'h17 : _GEN_1926; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1928 = 8'h88 == inBytes_7 ? 8'hc4 : _GEN_1927; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1929 = 8'h89 == inBytes_7 ? 8'ha7 : _GEN_1928; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1930 = 8'h8a == inBytes_7 ? 8'h7e : _GEN_1929; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1931 = 8'h8b == inBytes_7 ? 8'h3d : _GEN_1930; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1932 = 8'h8c == inBytes_7 ? 8'h64 : _GEN_1931; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1933 = 8'h8d == inBytes_7 ? 8'h5d : _GEN_1932; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1934 = 8'h8e == inBytes_7 ? 8'h19 : _GEN_1933; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1935 = 8'h8f == inBytes_7 ? 8'h73 : _GEN_1934; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1936 = 8'h90 == inBytes_7 ? 8'h60 : _GEN_1935; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1937 = 8'h91 == inBytes_7 ? 8'h81 : _GEN_1936; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1938 = 8'h92 == inBytes_7 ? 8'h4f : _GEN_1937; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1939 = 8'h93 == inBytes_7 ? 8'hdc : _GEN_1938; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1940 = 8'h94 == inBytes_7 ? 8'h22 : _GEN_1939; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1941 = 8'h95 == inBytes_7 ? 8'h2a : _GEN_1940; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1942 = 8'h96 == inBytes_7 ? 8'h90 : _GEN_1941; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1943 = 8'h97 == inBytes_7 ? 8'h88 : _GEN_1942; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1944 = 8'h98 == inBytes_7 ? 8'h46 : _GEN_1943; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1945 = 8'h99 == inBytes_7 ? 8'hee : _GEN_1944; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1946 = 8'h9a == inBytes_7 ? 8'hb8 : _GEN_1945; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1947 = 8'h9b == inBytes_7 ? 8'h14 : _GEN_1946; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1948 = 8'h9c == inBytes_7 ? 8'hde : _GEN_1947; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1949 = 8'h9d == inBytes_7 ? 8'h5e : _GEN_1948; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1950 = 8'h9e == inBytes_7 ? 8'hb : _GEN_1949; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1951 = 8'h9f == inBytes_7 ? 8'hdb : _GEN_1950; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1952 = 8'ha0 == inBytes_7 ? 8'he0 : _GEN_1951; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1953 = 8'ha1 == inBytes_7 ? 8'h32 : _GEN_1952; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1954 = 8'ha2 == inBytes_7 ? 8'h3a : _GEN_1953; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1955 = 8'ha3 == inBytes_7 ? 8'ha : _GEN_1954; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1956 = 8'ha4 == inBytes_7 ? 8'h49 : _GEN_1955; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1957 = 8'ha5 == inBytes_7 ? 8'h6 : _GEN_1956; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1958 = 8'ha6 == inBytes_7 ? 8'h24 : _GEN_1957; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1959 = 8'ha7 == inBytes_7 ? 8'h5c : _GEN_1958; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1960 = 8'ha8 == inBytes_7 ? 8'hc2 : _GEN_1959; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1961 = 8'ha9 == inBytes_7 ? 8'hd3 : _GEN_1960; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1962 = 8'haa == inBytes_7 ? 8'hac : _GEN_1961; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1963 = 8'hab == inBytes_7 ? 8'h62 : _GEN_1962; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1964 = 8'hac == inBytes_7 ? 8'h91 : _GEN_1963; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1965 = 8'had == inBytes_7 ? 8'h95 : _GEN_1964; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1966 = 8'hae == inBytes_7 ? 8'he4 : _GEN_1965; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1967 = 8'haf == inBytes_7 ? 8'h79 : _GEN_1966; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1968 = 8'hb0 == inBytes_7 ? 8'he7 : _GEN_1967; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1969 = 8'hb1 == inBytes_7 ? 8'hc8 : _GEN_1968; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1970 = 8'hb2 == inBytes_7 ? 8'h37 : _GEN_1969; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1971 = 8'hb3 == inBytes_7 ? 8'h6d : _GEN_1970; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1972 = 8'hb4 == inBytes_7 ? 8'h8d : _GEN_1971; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1973 = 8'hb5 == inBytes_7 ? 8'hd5 : _GEN_1972; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1974 = 8'hb6 == inBytes_7 ? 8'h4e : _GEN_1973; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1975 = 8'hb7 == inBytes_7 ? 8'ha9 : _GEN_1974; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1976 = 8'hb8 == inBytes_7 ? 8'h6c : _GEN_1975; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1977 = 8'hb9 == inBytes_7 ? 8'h56 : _GEN_1976; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1978 = 8'hba == inBytes_7 ? 8'hf4 : _GEN_1977; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1979 = 8'hbb == inBytes_7 ? 8'hea : _GEN_1978; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1980 = 8'hbc == inBytes_7 ? 8'h65 : _GEN_1979; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1981 = 8'hbd == inBytes_7 ? 8'h7a : _GEN_1980; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1982 = 8'hbe == inBytes_7 ? 8'hae : _GEN_1981; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1983 = 8'hbf == inBytes_7 ? 8'h8 : _GEN_1982; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1984 = 8'hc0 == inBytes_7 ? 8'hba : _GEN_1983; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1985 = 8'hc1 == inBytes_7 ? 8'h78 : _GEN_1984; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1986 = 8'hc2 == inBytes_7 ? 8'h25 : _GEN_1985; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1987 = 8'hc3 == inBytes_7 ? 8'h2e : _GEN_1986; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1988 = 8'hc4 == inBytes_7 ? 8'h1c : _GEN_1987; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1989 = 8'hc5 == inBytes_7 ? 8'ha6 : _GEN_1988; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1990 = 8'hc6 == inBytes_7 ? 8'hb4 : _GEN_1989; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1991 = 8'hc7 == inBytes_7 ? 8'hc6 : _GEN_1990; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1992 = 8'hc8 == inBytes_7 ? 8'he8 : _GEN_1991; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1993 = 8'hc9 == inBytes_7 ? 8'hdd : _GEN_1992; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1994 = 8'hca == inBytes_7 ? 8'h74 : _GEN_1993; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1995 = 8'hcb == inBytes_7 ? 8'h1f : _GEN_1994; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1996 = 8'hcc == inBytes_7 ? 8'h4b : _GEN_1995; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1997 = 8'hcd == inBytes_7 ? 8'hbd : _GEN_1996; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1998 = 8'hce == inBytes_7 ? 8'h8b : _GEN_1997; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_1999 = 8'hcf == inBytes_7 ? 8'h8a : _GEN_1998; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2000 = 8'hd0 == inBytes_7 ? 8'h70 : _GEN_1999; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2001 = 8'hd1 == inBytes_7 ? 8'h3e : _GEN_2000; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2002 = 8'hd2 == inBytes_7 ? 8'hb5 : _GEN_2001; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2003 = 8'hd3 == inBytes_7 ? 8'h66 : _GEN_2002; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2004 = 8'hd4 == inBytes_7 ? 8'h48 : _GEN_2003; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2005 = 8'hd5 == inBytes_7 ? 8'h3 : _GEN_2004; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2006 = 8'hd6 == inBytes_7 ? 8'hf6 : _GEN_2005; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2007 = 8'hd7 == inBytes_7 ? 8'he : _GEN_2006; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2008 = 8'hd8 == inBytes_7 ? 8'h61 : _GEN_2007; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2009 = 8'hd9 == inBytes_7 ? 8'h35 : _GEN_2008; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2010 = 8'hda == inBytes_7 ? 8'h57 : _GEN_2009; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2011 = 8'hdb == inBytes_7 ? 8'hb9 : _GEN_2010; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2012 = 8'hdc == inBytes_7 ? 8'h86 : _GEN_2011; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2013 = 8'hdd == inBytes_7 ? 8'hc1 : _GEN_2012; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2014 = 8'hde == inBytes_7 ? 8'h1d : _GEN_2013; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2015 = 8'hdf == inBytes_7 ? 8'h9e : _GEN_2014; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2016 = 8'he0 == inBytes_7 ? 8'he1 : _GEN_2015; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2017 = 8'he1 == inBytes_7 ? 8'hf8 : _GEN_2016; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2018 = 8'he2 == inBytes_7 ? 8'h98 : _GEN_2017; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2019 = 8'he3 == inBytes_7 ? 8'h11 : _GEN_2018; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2020 = 8'he4 == inBytes_7 ? 8'h69 : _GEN_2019; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2021 = 8'he5 == inBytes_7 ? 8'hd9 : _GEN_2020; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2022 = 8'he6 == inBytes_7 ? 8'h8e : _GEN_2021; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2023 = 8'he7 == inBytes_7 ? 8'h94 : _GEN_2022; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2024 = 8'he8 == inBytes_7 ? 8'h9b : _GEN_2023; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2025 = 8'he9 == inBytes_7 ? 8'h1e : _GEN_2024; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2026 = 8'hea == inBytes_7 ? 8'h87 : _GEN_2025; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2027 = 8'heb == inBytes_7 ? 8'he9 : _GEN_2026; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2028 = 8'hec == inBytes_7 ? 8'hce : _GEN_2027; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2029 = 8'hed == inBytes_7 ? 8'h55 : _GEN_2028; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2030 = 8'hee == inBytes_7 ? 8'h28 : _GEN_2029; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2031 = 8'hef == inBytes_7 ? 8'hdf : _GEN_2030; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2032 = 8'hf0 == inBytes_7 ? 8'h8c : _GEN_2031; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2033 = 8'hf1 == inBytes_7 ? 8'ha1 : _GEN_2032; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2034 = 8'hf2 == inBytes_7 ? 8'h89 : _GEN_2033; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2035 = 8'hf3 == inBytes_7 ? 8'hd : _GEN_2034; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2036 = 8'hf4 == inBytes_7 ? 8'hbf : _GEN_2035; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2037 = 8'hf5 == inBytes_7 ? 8'he6 : _GEN_2036; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2038 = 8'hf6 == inBytes_7 ? 8'h42 : _GEN_2037; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2039 = 8'hf7 == inBytes_7 ? 8'h68 : _GEN_2038; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2040 = 8'hf8 == inBytes_7 ? 8'h41 : _GEN_2039; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2041 = 8'hf9 == inBytes_7 ? 8'h99 : _GEN_2040; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2042 = 8'hfa == inBytes_7 ? 8'h2d : _GEN_2041; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2043 = 8'hfb == inBytes_7 ? 8'hf : _GEN_2042; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2044 = 8'hfc == inBytes_7 ? 8'hb0 : _GEN_2043; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2045 = 8'hfd == inBytes_7 ? 8'h54 : _GEN_2044; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2046 = 8'hfe == inBytes_7 ? 8'hbb : _GEN_2045; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] outBytes_7 = 8'hff == inBytes_7 ? 8'h16 : _GEN_2046; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2049 = 8'h1 == inBytes_8 ? 8'h7c : 8'h63; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2050 = 8'h2 == inBytes_8 ? 8'h77 : _GEN_2049; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2051 = 8'h3 == inBytes_8 ? 8'h7b : _GEN_2050; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2052 = 8'h4 == inBytes_8 ? 8'hf2 : _GEN_2051; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2053 = 8'h5 == inBytes_8 ? 8'h6b : _GEN_2052; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2054 = 8'h6 == inBytes_8 ? 8'h6f : _GEN_2053; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2055 = 8'h7 == inBytes_8 ? 8'hc5 : _GEN_2054; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2056 = 8'h8 == inBytes_8 ? 8'h30 : _GEN_2055; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2057 = 8'h9 == inBytes_8 ? 8'h1 : _GEN_2056; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2058 = 8'ha == inBytes_8 ? 8'h67 : _GEN_2057; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2059 = 8'hb == inBytes_8 ? 8'h2b : _GEN_2058; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2060 = 8'hc == inBytes_8 ? 8'hfe : _GEN_2059; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2061 = 8'hd == inBytes_8 ? 8'hd7 : _GEN_2060; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2062 = 8'he == inBytes_8 ? 8'hab : _GEN_2061; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2063 = 8'hf == inBytes_8 ? 8'h76 : _GEN_2062; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2064 = 8'h10 == inBytes_8 ? 8'hca : _GEN_2063; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2065 = 8'h11 == inBytes_8 ? 8'h82 : _GEN_2064; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2066 = 8'h12 == inBytes_8 ? 8'hc9 : _GEN_2065; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2067 = 8'h13 == inBytes_8 ? 8'h7d : _GEN_2066; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2068 = 8'h14 == inBytes_8 ? 8'hfa : _GEN_2067; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2069 = 8'h15 == inBytes_8 ? 8'h59 : _GEN_2068; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2070 = 8'h16 == inBytes_8 ? 8'h47 : _GEN_2069; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2071 = 8'h17 == inBytes_8 ? 8'hf0 : _GEN_2070; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2072 = 8'h18 == inBytes_8 ? 8'had : _GEN_2071; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2073 = 8'h19 == inBytes_8 ? 8'hd4 : _GEN_2072; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2074 = 8'h1a == inBytes_8 ? 8'ha2 : _GEN_2073; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2075 = 8'h1b == inBytes_8 ? 8'haf : _GEN_2074; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2076 = 8'h1c == inBytes_8 ? 8'h9c : _GEN_2075; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2077 = 8'h1d == inBytes_8 ? 8'ha4 : _GEN_2076; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2078 = 8'h1e == inBytes_8 ? 8'h72 : _GEN_2077; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2079 = 8'h1f == inBytes_8 ? 8'hc0 : _GEN_2078; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2080 = 8'h20 == inBytes_8 ? 8'hb7 : _GEN_2079; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2081 = 8'h21 == inBytes_8 ? 8'hfd : _GEN_2080; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2082 = 8'h22 == inBytes_8 ? 8'h93 : _GEN_2081; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2083 = 8'h23 == inBytes_8 ? 8'h26 : _GEN_2082; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2084 = 8'h24 == inBytes_8 ? 8'h36 : _GEN_2083; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2085 = 8'h25 == inBytes_8 ? 8'h3f : _GEN_2084; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2086 = 8'h26 == inBytes_8 ? 8'hf7 : _GEN_2085; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2087 = 8'h27 == inBytes_8 ? 8'hcc : _GEN_2086; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2088 = 8'h28 == inBytes_8 ? 8'h34 : _GEN_2087; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2089 = 8'h29 == inBytes_8 ? 8'ha5 : _GEN_2088; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2090 = 8'h2a == inBytes_8 ? 8'he5 : _GEN_2089; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2091 = 8'h2b == inBytes_8 ? 8'hf1 : _GEN_2090; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2092 = 8'h2c == inBytes_8 ? 8'h71 : _GEN_2091; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2093 = 8'h2d == inBytes_8 ? 8'hd8 : _GEN_2092; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2094 = 8'h2e == inBytes_8 ? 8'h31 : _GEN_2093; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2095 = 8'h2f == inBytes_8 ? 8'h15 : _GEN_2094; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2096 = 8'h30 == inBytes_8 ? 8'h4 : _GEN_2095; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2097 = 8'h31 == inBytes_8 ? 8'hc7 : _GEN_2096; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2098 = 8'h32 == inBytes_8 ? 8'h23 : _GEN_2097; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2099 = 8'h33 == inBytes_8 ? 8'hc3 : _GEN_2098; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2100 = 8'h34 == inBytes_8 ? 8'h18 : _GEN_2099; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2101 = 8'h35 == inBytes_8 ? 8'h96 : _GEN_2100; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2102 = 8'h36 == inBytes_8 ? 8'h5 : _GEN_2101; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2103 = 8'h37 == inBytes_8 ? 8'h9a : _GEN_2102; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2104 = 8'h38 == inBytes_8 ? 8'h7 : _GEN_2103; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2105 = 8'h39 == inBytes_8 ? 8'h12 : _GEN_2104; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2106 = 8'h3a == inBytes_8 ? 8'h80 : _GEN_2105; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2107 = 8'h3b == inBytes_8 ? 8'he2 : _GEN_2106; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2108 = 8'h3c == inBytes_8 ? 8'heb : _GEN_2107; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2109 = 8'h3d == inBytes_8 ? 8'h27 : _GEN_2108; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2110 = 8'h3e == inBytes_8 ? 8'hb2 : _GEN_2109; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2111 = 8'h3f == inBytes_8 ? 8'h75 : _GEN_2110; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2112 = 8'h40 == inBytes_8 ? 8'h9 : _GEN_2111; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2113 = 8'h41 == inBytes_8 ? 8'h83 : _GEN_2112; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2114 = 8'h42 == inBytes_8 ? 8'h2c : _GEN_2113; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2115 = 8'h43 == inBytes_8 ? 8'h1a : _GEN_2114; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2116 = 8'h44 == inBytes_8 ? 8'h1b : _GEN_2115; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2117 = 8'h45 == inBytes_8 ? 8'h6e : _GEN_2116; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2118 = 8'h46 == inBytes_8 ? 8'h5a : _GEN_2117; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2119 = 8'h47 == inBytes_8 ? 8'ha0 : _GEN_2118; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2120 = 8'h48 == inBytes_8 ? 8'h52 : _GEN_2119; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2121 = 8'h49 == inBytes_8 ? 8'h3b : _GEN_2120; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2122 = 8'h4a == inBytes_8 ? 8'hd6 : _GEN_2121; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2123 = 8'h4b == inBytes_8 ? 8'hb3 : _GEN_2122; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2124 = 8'h4c == inBytes_8 ? 8'h29 : _GEN_2123; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2125 = 8'h4d == inBytes_8 ? 8'he3 : _GEN_2124; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2126 = 8'h4e == inBytes_8 ? 8'h2f : _GEN_2125; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2127 = 8'h4f == inBytes_8 ? 8'h84 : _GEN_2126; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2128 = 8'h50 == inBytes_8 ? 8'h53 : _GEN_2127; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2129 = 8'h51 == inBytes_8 ? 8'hd1 : _GEN_2128; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2130 = 8'h52 == inBytes_8 ? 8'h0 : _GEN_2129; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2131 = 8'h53 == inBytes_8 ? 8'hed : _GEN_2130; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2132 = 8'h54 == inBytes_8 ? 8'h20 : _GEN_2131; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2133 = 8'h55 == inBytes_8 ? 8'hfc : _GEN_2132; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2134 = 8'h56 == inBytes_8 ? 8'hb1 : _GEN_2133; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2135 = 8'h57 == inBytes_8 ? 8'h5b : _GEN_2134; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2136 = 8'h58 == inBytes_8 ? 8'h6a : _GEN_2135; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2137 = 8'h59 == inBytes_8 ? 8'hcb : _GEN_2136; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2138 = 8'h5a == inBytes_8 ? 8'hbe : _GEN_2137; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2139 = 8'h5b == inBytes_8 ? 8'h39 : _GEN_2138; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2140 = 8'h5c == inBytes_8 ? 8'h4a : _GEN_2139; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2141 = 8'h5d == inBytes_8 ? 8'h4c : _GEN_2140; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2142 = 8'h5e == inBytes_8 ? 8'h58 : _GEN_2141; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2143 = 8'h5f == inBytes_8 ? 8'hcf : _GEN_2142; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2144 = 8'h60 == inBytes_8 ? 8'hd0 : _GEN_2143; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2145 = 8'h61 == inBytes_8 ? 8'hef : _GEN_2144; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2146 = 8'h62 == inBytes_8 ? 8'haa : _GEN_2145; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2147 = 8'h63 == inBytes_8 ? 8'hfb : _GEN_2146; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2148 = 8'h64 == inBytes_8 ? 8'h43 : _GEN_2147; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2149 = 8'h65 == inBytes_8 ? 8'h4d : _GEN_2148; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2150 = 8'h66 == inBytes_8 ? 8'h33 : _GEN_2149; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2151 = 8'h67 == inBytes_8 ? 8'h85 : _GEN_2150; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2152 = 8'h68 == inBytes_8 ? 8'h45 : _GEN_2151; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2153 = 8'h69 == inBytes_8 ? 8'hf9 : _GEN_2152; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2154 = 8'h6a == inBytes_8 ? 8'h2 : _GEN_2153; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2155 = 8'h6b == inBytes_8 ? 8'h7f : _GEN_2154; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2156 = 8'h6c == inBytes_8 ? 8'h50 : _GEN_2155; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2157 = 8'h6d == inBytes_8 ? 8'h3c : _GEN_2156; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2158 = 8'h6e == inBytes_8 ? 8'h9f : _GEN_2157; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2159 = 8'h6f == inBytes_8 ? 8'ha8 : _GEN_2158; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2160 = 8'h70 == inBytes_8 ? 8'h51 : _GEN_2159; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2161 = 8'h71 == inBytes_8 ? 8'ha3 : _GEN_2160; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2162 = 8'h72 == inBytes_8 ? 8'h40 : _GEN_2161; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2163 = 8'h73 == inBytes_8 ? 8'h8f : _GEN_2162; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2164 = 8'h74 == inBytes_8 ? 8'h92 : _GEN_2163; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2165 = 8'h75 == inBytes_8 ? 8'h9d : _GEN_2164; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2166 = 8'h76 == inBytes_8 ? 8'h38 : _GEN_2165; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2167 = 8'h77 == inBytes_8 ? 8'hf5 : _GEN_2166; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2168 = 8'h78 == inBytes_8 ? 8'hbc : _GEN_2167; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2169 = 8'h79 == inBytes_8 ? 8'hb6 : _GEN_2168; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2170 = 8'h7a == inBytes_8 ? 8'hda : _GEN_2169; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2171 = 8'h7b == inBytes_8 ? 8'h21 : _GEN_2170; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2172 = 8'h7c == inBytes_8 ? 8'h10 : _GEN_2171; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2173 = 8'h7d == inBytes_8 ? 8'hff : _GEN_2172; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2174 = 8'h7e == inBytes_8 ? 8'hf3 : _GEN_2173; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2175 = 8'h7f == inBytes_8 ? 8'hd2 : _GEN_2174; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2176 = 8'h80 == inBytes_8 ? 8'hcd : _GEN_2175; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2177 = 8'h81 == inBytes_8 ? 8'hc : _GEN_2176; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2178 = 8'h82 == inBytes_8 ? 8'h13 : _GEN_2177; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2179 = 8'h83 == inBytes_8 ? 8'hec : _GEN_2178; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2180 = 8'h84 == inBytes_8 ? 8'h5f : _GEN_2179; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2181 = 8'h85 == inBytes_8 ? 8'h97 : _GEN_2180; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2182 = 8'h86 == inBytes_8 ? 8'h44 : _GEN_2181; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2183 = 8'h87 == inBytes_8 ? 8'h17 : _GEN_2182; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2184 = 8'h88 == inBytes_8 ? 8'hc4 : _GEN_2183; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2185 = 8'h89 == inBytes_8 ? 8'ha7 : _GEN_2184; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2186 = 8'h8a == inBytes_8 ? 8'h7e : _GEN_2185; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2187 = 8'h8b == inBytes_8 ? 8'h3d : _GEN_2186; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2188 = 8'h8c == inBytes_8 ? 8'h64 : _GEN_2187; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2189 = 8'h8d == inBytes_8 ? 8'h5d : _GEN_2188; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2190 = 8'h8e == inBytes_8 ? 8'h19 : _GEN_2189; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2191 = 8'h8f == inBytes_8 ? 8'h73 : _GEN_2190; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2192 = 8'h90 == inBytes_8 ? 8'h60 : _GEN_2191; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2193 = 8'h91 == inBytes_8 ? 8'h81 : _GEN_2192; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2194 = 8'h92 == inBytes_8 ? 8'h4f : _GEN_2193; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2195 = 8'h93 == inBytes_8 ? 8'hdc : _GEN_2194; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2196 = 8'h94 == inBytes_8 ? 8'h22 : _GEN_2195; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2197 = 8'h95 == inBytes_8 ? 8'h2a : _GEN_2196; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2198 = 8'h96 == inBytes_8 ? 8'h90 : _GEN_2197; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2199 = 8'h97 == inBytes_8 ? 8'h88 : _GEN_2198; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2200 = 8'h98 == inBytes_8 ? 8'h46 : _GEN_2199; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2201 = 8'h99 == inBytes_8 ? 8'hee : _GEN_2200; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2202 = 8'h9a == inBytes_8 ? 8'hb8 : _GEN_2201; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2203 = 8'h9b == inBytes_8 ? 8'h14 : _GEN_2202; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2204 = 8'h9c == inBytes_8 ? 8'hde : _GEN_2203; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2205 = 8'h9d == inBytes_8 ? 8'h5e : _GEN_2204; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2206 = 8'h9e == inBytes_8 ? 8'hb : _GEN_2205; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2207 = 8'h9f == inBytes_8 ? 8'hdb : _GEN_2206; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2208 = 8'ha0 == inBytes_8 ? 8'he0 : _GEN_2207; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2209 = 8'ha1 == inBytes_8 ? 8'h32 : _GEN_2208; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2210 = 8'ha2 == inBytes_8 ? 8'h3a : _GEN_2209; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2211 = 8'ha3 == inBytes_8 ? 8'ha : _GEN_2210; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2212 = 8'ha4 == inBytes_8 ? 8'h49 : _GEN_2211; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2213 = 8'ha5 == inBytes_8 ? 8'h6 : _GEN_2212; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2214 = 8'ha6 == inBytes_8 ? 8'h24 : _GEN_2213; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2215 = 8'ha7 == inBytes_8 ? 8'h5c : _GEN_2214; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2216 = 8'ha8 == inBytes_8 ? 8'hc2 : _GEN_2215; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2217 = 8'ha9 == inBytes_8 ? 8'hd3 : _GEN_2216; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2218 = 8'haa == inBytes_8 ? 8'hac : _GEN_2217; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2219 = 8'hab == inBytes_8 ? 8'h62 : _GEN_2218; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2220 = 8'hac == inBytes_8 ? 8'h91 : _GEN_2219; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2221 = 8'had == inBytes_8 ? 8'h95 : _GEN_2220; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2222 = 8'hae == inBytes_8 ? 8'he4 : _GEN_2221; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2223 = 8'haf == inBytes_8 ? 8'h79 : _GEN_2222; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2224 = 8'hb0 == inBytes_8 ? 8'he7 : _GEN_2223; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2225 = 8'hb1 == inBytes_8 ? 8'hc8 : _GEN_2224; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2226 = 8'hb2 == inBytes_8 ? 8'h37 : _GEN_2225; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2227 = 8'hb3 == inBytes_8 ? 8'h6d : _GEN_2226; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2228 = 8'hb4 == inBytes_8 ? 8'h8d : _GEN_2227; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2229 = 8'hb5 == inBytes_8 ? 8'hd5 : _GEN_2228; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2230 = 8'hb6 == inBytes_8 ? 8'h4e : _GEN_2229; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2231 = 8'hb7 == inBytes_8 ? 8'ha9 : _GEN_2230; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2232 = 8'hb8 == inBytes_8 ? 8'h6c : _GEN_2231; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2233 = 8'hb9 == inBytes_8 ? 8'h56 : _GEN_2232; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2234 = 8'hba == inBytes_8 ? 8'hf4 : _GEN_2233; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2235 = 8'hbb == inBytes_8 ? 8'hea : _GEN_2234; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2236 = 8'hbc == inBytes_8 ? 8'h65 : _GEN_2235; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2237 = 8'hbd == inBytes_8 ? 8'h7a : _GEN_2236; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2238 = 8'hbe == inBytes_8 ? 8'hae : _GEN_2237; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2239 = 8'hbf == inBytes_8 ? 8'h8 : _GEN_2238; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2240 = 8'hc0 == inBytes_8 ? 8'hba : _GEN_2239; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2241 = 8'hc1 == inBytes_8 ? 8'h78 : _GEN_2240; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2242 = 8'hc2 == inBytes_8 ? 8'h25 : _GEN_2241; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2243 = 8'hc3 == inBytes_8 ? 8'h2e : _GEN_2242; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2244 = 8'hc4 == inBytes_8 ? 8'h1c : _GEN_2243; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2245 = 8'hc5 == inBytes_8 ? 8'ha6 : _GEN_2244; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2246 = 8'hc6 == inBytes_8 ? 8'hb4 : _GEN_2245; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2247 = 8'hc7 == inBytes_8 ? 8'hc6 : _GEN_2246; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2248 = 8'hc8 == inBytes_8 ? 8'he8 : _GEN_2247; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2249 = 8'hc9 == inBytes_8 ? 8'hdd : _GEN_2248; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2250 = 8'hca == inBytes_8 ? 8'h74 : _GEN_2249; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2251 = 8'hcb == inBytes_8 ? 8'h1f : _GEN_2250; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2252 = 8'hcc == inBytes_8 ? 8'h4b : _GEN_2251; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2253 = 8'hcd == inBytes_8 ? 8'hbd : _GEN_2252; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2254 = 8'hce == inBytes_8 ? 8'h8b : _GEN_2253; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2255 = 8'hcf == inBytes_8 ? 8'h8a : _GEN_2254; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2256 = 8'hd0 == inBytes_8 ? 8'h70 : _GEN_2255; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2257 = 8'hd1 == inBytes_8 ? 8'h3e : _GEN_2256; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2258 = 8'hd2 == inBytes_8 ? 8'hb5 : _GEN_2257; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2259 = 8'hd3 == inBytes_8 ? 8'h66 : _GEN_2258; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2260 = 8'hd4 == inBytes_8 ? 8'h48 : _GEN_2259; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2261 = 8'hd5 == inBytes_8 ? 8'h3 : _GEN_2260; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2262 = 8'hd6 == inBytes_8 ? 8'hf6 : _GEN_2261; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2263 = 8'hd7 == inBytes_8 ? 8'he : _GEN_2262; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2264 = 8'hd8 == inBytes_8 ? 8'h61 : _GEN_2263; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2265 = 8'hd9 == inBytes_8 ? 8'h35 : _GEN_2264; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2266 = 8'hda == inBytes_8 ? 8'h57 : _GEN_2265; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2267 = 8'hdb == inBytes_8 ? 8'hb9 : _GEN_2266; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2268 = 8'hdc == inBytes_8 ? 8'h86 : _GEN_2267; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2269 = 8'hdd == inBytes_8 ? 8'hc1 : _GEN_2268; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2270 = 8'hde == inBytes_8 ? 8'h1d : _GEN_2269; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2271 = 8'hdf == inBytes_8 ? 8'h9e : _GEN_2270; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2272 = 8'he0 == inBytes_8 ? 8'he1 : _GEN_2271; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2273 = 8'he1 == inBytes_8 ? 8'hf8 : _GEN_2272; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2274 = 8'he2 == inBytes_8 ? 8'h98 : _GEN_2273; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2275 = 8'he3 == inBytes_8 ? 8'h11 : _GEN_2274; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2276 = 8'he4 == inBytes_8 ? 8'h69 : _GEN_2275; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2277 = 8'he5 == inBytes_8 ? 8'hd9 : _GEN_2276; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2278 = 8'he6 == inBytes_8 ? 8'h8e : _GEN_2277; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2279 = 8'he7 == inBytes_8 ? 8'h94 : _GEN_2278; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2280 = 8'he8 == inBytes_8 ? 8'h9b : _GEN_2279; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2281 = 8'he9 == inBytes_8 ? 8'h1e : _GEN_2280; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2282 = 8'hea == inBytes_8 ? 8'h87 : _GEN_2281; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2283 = 8'heb == inBytes_8 ? 8'he9 : _GEN_2282; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2284 = 8'hec == inBytes_8 ? 8'hce : _GEN_2283; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2285 = 8'hed == inBytes_8 ? 8'h55 : _GEN_2284; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2286 = 8'hee == inBytes_8 ? 8'h28 : _GEN_2285; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2287 = 8'hef == inBytes_8 ? 8'hdf : _GEN_2286; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2288 = 8'hf0 == inBytes_8 ? 8'h8c : _GEN_2287; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2289 = 8'hf1 == inBytes_8 ? 8'ha1 : _GEN_2288; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2290 = 8'hf2 == inBytes_8 ? 8'h89 : _GEN_2289; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2291 = 8'hf3 == inBytes_8 ? 8'hd : _GEN_2290; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2292 = 8'hf4 == inBytes_8 ? 8'hbf : _GEN_2291; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2293 = 8'hf5 == inBytes_8 ? 8'he6 : _GEN_2292; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2294 = 8'hf6 == inBytes_8 ? 8'h42 : _GEN_2293; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2295 = 8'hf7 == inBytes_8 ? 8'h68 : _GEN_2294; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2296 = 8'hf8 == inBytes_8 ? 8'h41 : _GEN_2295; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2297 = 8'hf9 == inBytes_8 ? 8'h99 : _GEN_2296; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2298 = 8'hfa == inBytes_8 ? 8'h2d : _GEN_2297; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2299 = 8'hfb == inBytes_8 ? 8'hf : _GEN_2298; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2300 = 8'hfc == inBytes_8 ? 8'hb0 : _GEN_2299; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2301 = 8'hfd == inBytes_8 ? 8'h54 : _GEN_2300; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2302 = 8'hfe == inBytes_8 ? 8'hbb : _GEN_2301; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] outBytes_8 = 8'hff == inBytes_8 ? 8'h16 : _GEN_2302; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2305 = 8'h1 == inBytes_9 ? 8'h7c : 8'h63; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2306 = 8'h2 == inBytes_9 ? 8'h77 : _GEN_2305; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2307 = 8'h3 == inBytes_9 ? 8'h7b : _GEN_2306; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2308 = 8'h4 == inBytes_9 ? 8'hf2 : _GEN_2307; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2309 = 8'h5 == inBytes_9 ? 8'h6b : _GEN_2308; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2310 = 8'h6 == inBytes_9 ? 8'h6f : _GEN_2309; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2311 = 8'h7 == inBytes_9 ? 8'hc5 : _GEN_2310; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2312 = 8'h8 == inBytes_9 ? 8'h30 : _GEN_2311; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2313 = 8'h9 == inBytes_9 ? 8'h1 : _GEN_2312; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2314 = 8'ha == inBytes_9 ? 8'h67 : _GEN_2313; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2315 = 8'hb == inBytes_9 ? 8'h2b : _GEN_2314; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2316 = 8'hc == inBytes_9 ? 8'hfe : _GEN_2315; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2317 = 8'hd == inBytes_9 ? 8'hd7 : _GEN_2316; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2318 = 8'he == inBytes_9 ? 8'hab : _GEN_2317; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2319 = 8'hf == inBytes_9 ? 8'h76 : _GEN_2318; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2320 = 8'h10 == inBytes_9 ? 8'hca : _GEN_2319; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2321 = 8'h11 == inBytes_9 ? 8'h82 : _GEN_2320; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2322 = 8'h12 == inBytes_9 ? 8'hc9 : _GEN_2321; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2323 = 8'h13 == inBytes_9 ? 8'h7d : _GEN_2322; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2324 = 8'h14 == inBytes_9 ? 8'hfa : _GEN_2323; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2325 = 8'h15 == inBytes_9 ? 8'h59 : _GEN_2324; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2326 = 8'h16 == inBytes_9 ? 8'h47 : _GEN_2325; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2327 = 8'h17 == inBytes_9 ? 8'hf0 : _GEN_2326; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2328 = 8'h18 == inBytes_9 ? 8'had : _GEN_2327; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2329 = 8'h19 == inBytes_9 ? 8'hd4 : _GEN_2328; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2330 = 8'h1a == inBytes_9 ? 8'ha2 : _GEN_2329; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2331 = 8'h1b == inBytes_9 ? 8'haf : _GEN_2330; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2332 = 8'h1c == inBytes_9 ? 8'h9c : _GEN_2331; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2333 = 8'h1d == inBytes_9 ? 8'ha4 : _GEN_2332; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2334 = 8'h1e == inBytes_9 ? 8'h72 : _GEN_2333; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2335 = 8'h1f == inBytes_9 ? 8'hc0 : _GEN_2334; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2336 = 8'h20 == inBytes_9 ? 8'hb7 : _GEN_2335; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2337 = 8'h21 == inBytes_9 ? 8'hfd : _GEN_2336; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2338 = 8'h22 == inBytes_9 ? 8'h93 : _GEN_2337; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2339 = 8'h23 == inBytes_9 ? 8'h26 : _GEN_2338; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2340 = 8'h24 == inBytes_9 ? 8'h36 : _GEN_2339; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2341 = 8'h25 == inBytes_9 ? 8'h3f : _GEN_2340; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2342 = 8'h26 == inBytes_9 ? 8'hf7 : _GEN_2341; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2343 = 8'h27 == inBytes_9 ? 8'hcc : _GEN_2342; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2344 = 8'h28 == inBytes_9 ? 8'h34 : _GEN_2343; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2345 = 8'h29 == inBytes_9 ? 8'ha5 : _GEN_2344; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2346 = 8'h2a == inBytes_9 ? 8'he5 : _GEN_2345; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2347 = 8'h2b == inBytes_9 ? 8'hf1 : _GEN_2346; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2348 = 8'h2c == inBytes_9 ? 8'h71 : _GEN_2347; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2349 = 8'h2d == inBytes_9 ? 8'hd8 : _GEN_2348; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2350 = 8'h2e == inBytes_9 ? 8'h31 : _GEN_2349; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2351 = 8'h2f == inBytes_9 ? 8'h15 : _GEN_2350; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2352 = 8'h30 == inBytes_9 ? 8'h4 : _GEN_2351; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2353 = 8'h31 == inBytes_9 ? 8'hc7 : _GEN_2352; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2354 = 8'h32 == inBytes_9 ? 8'h23 : _GEN_2353; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2355 = 8'h33 == inBytes_9 ? 8'hc3 : _GEN_2354; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2356 = 8'h34 == inBytes_9 ? 8'h18 : _GEN_2355; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2357 = 8'h35 == inBytes_9 ? 8'h96 : _GEN_2356; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2358 = 8'h36 == inBytes_9 ? 8'h5 : _GEN_2357; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2359 = 8'h37 == inBytes_9 ? 8'h9a : _GEN_2358; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2360 = 8'h38 == inBytes_9 ? 8'h7 : _GEN_2359; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2361 = 8'h39 == inBytes_9 ? 8'h12 : _GEN_2360; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2362 = 8'h3a == inBytes_9 ? 8'h80 : _GEN_2361; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2363 = 8'h3b == inBytes_9 ? 8'he2 : _GEN_2362; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2364 = 8'h3c == inBytes_9 ? 8'heb : _GEN_2363; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2365 = 8'h3d == inBytes_9 ? 8'h27 : _GEN_2364; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2366 = 8'h3e == inBytes_9 ? 8'hb2 : _GEN_2365; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2367 = 8'h3f == inBytes_9 ? 8'h75 : _GEN_2366; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2368 = 8'h40 == inBytes_9 ? 8'h9 : _GEN_2367; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2369 = 8'h41 == inBytes_9 ? 8'h83 : _GEN_2368; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2370 = 8'h42 == inBytes_9 ? 8'h2c : _GEN_2369; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2371 = 8'h43 == inBytes_9 ? 8'h1a : _GEN_2370; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2372 = 8'h44 == inBytes_9 ? 8'h1b : _GEN_2371; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2373 = 8'h45 == inBytes_9 ? 8'h6e : _GEN_2372; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2374 = 8'h46 == inBytes_9 ? 8'h5a : _GEN_2373; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2375 = 8'h47 == inBytes_9 ? 8'ha0 : _GEN_2374; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2376 = 8'h48 == inBytes_9 ? 8'h52 : _GEN_2375; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2377 = 8'h49 == inBytes_9 ? 8'h3b : _GEN_2376; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2378 = 8'h4a == inBytes_9 ? 8'hd6 : _GEN_2377; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2379 = 8'h4b == inBytes_9 ? 8'hb3 : _GEN_2378; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2380 = 8'h4c == inBytes_9 ? 8'h29 : _GEN_2379; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2381 = 8'h4d == inBytes_9 ? 8'he3 : _GEN_2380; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2382 = 8'h4e == inBytes_9 ? 8'h2f : _GEN_2381; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2383 = 8'h4f == inBytes_9 ? 8'h84 : _GEN_2382; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2384 = 8'h50 == inBytes_9 ? 8'h53 : _GEN_2383; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2385 = 8'h51 == inBytes_9 ? 8'hd1 : _GEN_2384; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2386 = 8'h52 == inBytes_9 ? 8'h0 : _GEN_2385; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2387 = 8'h53 == inBytes_9 ? 8'hed : _GEN_2386; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2388 = 8'h54 == inBytes_9 ? 8'h20 : _GEN_2387; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2389 = 8'h55 == inBytes_9 ? 8'hfc : _GEN_2388; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2390 = 8'h56 == inBytes_9 ? 8'hb1 : _GEN_2389; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2391 = 8'h57 == inBytes_9 ? 8'h5b : _GEN_2390; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2392 = 8'h58 == inBytes_9 ? 8'h6a : _GEN_2391; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2393 = 8'h59 == inBytes_9 ? 8'hcb : _GEN_2392; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2394 = 8'h5a == inBytes_9 ? 8'hbe : _GEN_2393; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2395 = 8'h5b == inBytes_9 ? 8'h39 : _GEN_2394; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2396 = 8'h5c == inBytes_9 ? 8'h4a : _GEN_2395; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2397 = 8'h5d == inBytes_9 ? 8'h4c : _GEN_2396; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2398 = 8'h5e == inBytes_9 ? 8'h58 : _GEN_2397; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2399 = 8'h5f == inBytes_9 ? 8'hcf : _GEN_2398; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2400 = 8'h60 == inBytes_9 ? 8'hd0 : _GEN_2399; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2401 = 8'h61 == inBytes_9 ? 8'hef : _GEN_2400; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2402 = 8'h62 == inBytes_9 ? 8'haa : _GEN_2401; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2403 = 8'h63 == inBytes_9 ? 8'hfb : _GEN_2402; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2404 = 8'h64 == inBytes_9 ? 8'h43 : _GEN_2403; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2405 = 8'h65 == inBytes_9 ? 8'h4d : _GEN_2404; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2406 = 8'h66 == inBytes_9 ? 8'h33 : _GEN_2405; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2407 = 8'h67 == inBytes_9 ? 8'h85 : _GEN_2406; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2408 = 8'h68 == inBytes_9 ? 8'h45 : _GEN_2407; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2409 = 8'h69 == inBytes_9 ? 8'hf9 : _GEN_2408; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2410 = 8'h6a == inBytes_9 ? 8'h2 : _GEN_2409; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2411 = 8'h6b == inBytes_9 ? 8'h7f : _GEN_2410; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2412 = 8'h6c == inBytes_9 ? 8'h50 : _GEN_2411; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2413 = 8'h6d == inBytes_9 ? 8'h3c : _GEN_2412; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2414 = 8'h6e == inBytes_9 ? 8'h9f : _GEN_2413; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2415 = 8'h6f == inBytes_9 ? 8'ha8 : _GEN_2414; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2416 = 8'h70 == inBytes_9 ? 8'h51 : _GEN_2415; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2417 = 8'h71 == inBytes_9 ? 8'ha3 : _GEN_2416; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2418 = 8'h72 == inBytes_9 ? 8'h40 : _GEN_2417; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2419 = 8'h73 == inBytes_9 ? 8'h8f : _GEN_2418; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2420 = 8'h74 == inBytes_9 ? 8'h92 : _GEN_2419; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2421 = 8'h75 == inBytes_9 ? 8'h9d : _GEN_2420; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2422 = 8'h76 == inBytes_9 ? 8'h38 : _GEN_2421; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2423 = 8'h77 == inBytes_9 ? 8'hf5 : _GEN_2422; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2424 = 8'h78 == inBytes_9 ? 8'hbc : _GEN_2423; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2425 = 8'h79 == inBytes_9 ? 8'hb6 : _GEN_2424; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2426 = 8'h7a == inBytes_9 ? 8'hda : _GEN_2425; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2427 = 8'h7b == inBytes_9 ? 8'h21 : _GEN_2426; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2428 = 8'h7c == inBytes_9 ? 8'h10 : _GEN_2427; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2429 = 8'h7d == inBytes_9 ? 8'hff : _GEN_2428; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2430 = 8'h7e == inBytes_9 ? 8'hf3 : _GEN_2429; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2431 = 8'h7f == inBytes_9 ? 8'hd2 : _GEN_2430; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2432 = 8'h80 == inBytes_9 ? 8'hcd : _GEN_2431; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2433 = 8'h81 == inBytes_9 ? 8'hc : _GEN_2432; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2434 = 8'h82 == inBytes_9 ? 8'h13 : _GEN_2433; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2435 = 8'h83 == inBytes_9 ? 8'hec : _GEN_2434; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2436 = 8'h84 == inBytes_9 ? 8'h5f : _GEN_2435; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2437 = 8'h85 == inBytes_9 ? 8'h97 : _GEN_2436; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2438 = 8'h86 == inBytes_9 ? 8'h44 : _GEN_2437; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2439 = 8'h87 == inBytes_9 ? 8'h17 : _GEN_2438; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2440 = 8'h88 == inBytes_9 ? 8'hc4 : _GEN_2439; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2441 = 8'h89 == inBytes_9 ? 8'ha7 : _GEN_2440; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2442 = 8'h8a == inBytes_9 ? 8'h7e : _GEN_2441; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2443 = 8'h8b == inBytes_9 ? 8'h3d : _GEN_2442; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2444 = 8'h8c == inBytes_9 ? 8'h64 : _GEN_2443; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2445 = 8'h8d == inBytes_9 ? 8'h5d : _GEN_2444; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2446 = 8'h8e == inBytes_9 ? 8'h19 : _GEN_2445; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2447 = 8'h8f == inBytes_9 ? 8'h73 : _GEN_2446; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2448 = 8'h90 == inBytes_9 ? 8'h60 : _GEN_2447; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2449 = 8'h91 == inBytes_9 ? 8'h81 : _GEN_2448; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2450 = 8'h92 == inBytes_9 ? 8'h4f : _GEN_2449; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2451 = 8'h93 == inBytes_9 ? 8'hdc : _GEN_2450; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2452 = 8'h94 == inBytes_9 ? 8'h22 : _GEN_2451; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2453 = 8'h95 == inBytes_9 ? 8'h2a : _GEN_2452; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2454 = 8'h96 == inBytes_9 ? 8'h90 : _GEN_2453; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2455 = 8'h97 == inBytes_9 ? 8'h88 : _GEN_2454; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2456 = 8'h98 == inBytes_9 ? 8'h46 : _GEN_2455; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2457 = 8'h99 == inBytes_9 ? 8'hee : _GEN_2456; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2458 = 8'h9a == inBytes_9 ? 8'hb8 : _GEN_2457; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2459 = 8'h9b == inBytes_9 ? 8'h14 : _GEN_2458; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2460 = 8'h9c == inBytes_9 ? 8'hde : _GEN_2459; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2461 = 8'h9d == inBytes_9 ? 8'h5e : _GEN_2460; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2462 = 8'h9e == inBytes_9 ? 8'hb : _GEN_2461; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2463 = 8'h9f == inBytes_9 ? 8'hdb : _GEN_2462; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2464 = 8'ha0 == inBytes_9 ? 8'he0 : _GEN_2463; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2465 = 8'ha1 == inBytes_9 ? 8'h32 : _GEN_2464; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2466 = 8'ha2 == inBytes_9 ? 8'h3a : _GEN_2465; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2467 = 8'ha3 == inBytes_9 ? 8'ha : _GEN_2466; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2468 = 8'ha4 == inBytes_9 ? 8'h49 : _GEN_2467; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2469 = 8'ha5 == inBytes_9 ? 8'h6 : _GEN_2468; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2470 = 8'ha6 == inBytes_9 ? 8'h24 : _GEN_2469; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2471 = 8'ha7 == inBytes_9 ? 8'h5c : _GEN_2470; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2472 = 8'ha8 == inBytes_9 ? 8'hc2 : _GEN_2471; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2473 = 8'ha9 == inBytes_9 ? 8'hd3 : _GEN_2472; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2474 = 8'haa == inBytes_9 ? 8'hac : _GEN_2473; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2475 = 8'hab == inBytes_9 ? 8'h62 : _GEN_2474; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2476 = 8'hac == inBytes_9 ? 8'h91 : _GEN_2475; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2477 = 8'had == inBytes_9 ? 8'h95 : _GEN_2476; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2478 = 8'hae == inBytes_9 ? 8'he4 : _GEN_2477; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2479 = 8'haf == inBytes_9 ? 8'h79 : _GEN_2478; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2480 = 8'hb0 == inBytes_9 ? 8'he7 : _GEN_2479; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2481 = 8'hb1 == inBytes_9 ? 8'hc8 : _GEN_2480; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2482 = 8'hb2 == inBytes_9 ? 8'h37 : _GEN_2481; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2483 = 8'hb3 == inBytes_9 ? 8'h6d : _GEN_2482; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2484 = 8'hb4 == inBytes_9 ? 8'h8d : _GEN_2483; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2485 = 8'hb5 == inBytes_9 ? 8'hd5 : _GEN_2484; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2486 = 8'hb6 == inBytes_9 ? 8'h4e : _GEN_2485; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2487 = 8'hb7 == inBytes_9 ? 8'ha9 : _GEN_2486; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2488 = 8'hb8 == inBytes_9 ? 8'h6c : _GEN_2487; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2489 = 8'hb9 == inBytes_9 ? 8'h56 : _GEN_2488; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2490 = 8'hba == inBytes_9 ? 8'hf4 : _GEN_2489; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2491 = 8'hbb == inBytes_9 ? 8'hea : _GEN_2490; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2492 = 8'hbc == inBytes_9 ? 8'h65 : _GEN_2491; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2493 = 8'hbd == inBytes_9 ? 8'h7a : _GEN_2492; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2494 = 8'hbe == inBytes_9 ? 8'hae : _GEN_2493; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2495 = 8'hbf == inBytes_9 ? 8'h8 : _GEN_2494; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2496 = 8'hc0 == inBytes_9 ? 8'hba : _GEN_2495; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2497 = 8'hc1 == inBytes_9 ? 8'h78 : _GEN_2496; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2498 = 8'hc2 == inBytes_9 ? 8'h25 : _GEN_2497; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2499 = 8'hc3 == inBytes_9 ? 8'h2e : _GEN_2498; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2500 = 8'hc4 == inBytes_9 ? 8'h1c : _GEN_2499; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2501 = 8'hc5 == inBytes_9 ? 8'ha6 : _GEN_2500; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2502 = 8'hc6 == inBytes_9 ? 8'hb4 : _GEN_2501; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2503 = 8'hc7 == inBytes_9 ? 8'hc6 : _GEN_2502; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2504 = 8'hc8 == inBytes_9 ? 8'he8 : _GEN_2503; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2505 = 8'hc9 == inBytes_9 ? 8'hdd : _GEN_2504; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2506 = 8'hca == inBytes_9 ? 8'h74 : _GEN_2505; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2507 = 8'hcb == inBytes_9 ? 8'h1f : _GEN_2506; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2508 = 8'hcc == inBytes_9 ? 8'h4b : _GEN_2507; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2509 = 8'hcd == inBytes_9 ? 8'hbd : _GEN_2508; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2510 = 8'hce == inBytes_9 ? 8'h8b : _GEN_2509; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2511 = 8'hcf == inBytes_9 ? 8'h8a : _GEN_2510; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2512 = 8'hd0 == inBytes_9 ? 8'h70 : _GEN_2511; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2513 = 8'hd1 == inBytes_9 ? 8'h3e : _GEN_2512; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2514 = 8'hd2 == inBytes_9 ? 8'hb5 : _GEN_2513; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2515 = 8'hd3 == inBytes_9 ? 8'h66 : _GEN_2514; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2516 = 8'hd4 == inBytes_9 ? 8'h48 : _GEN_2515; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2517 = 8'hd5 == inBytes_9 ? 8'h3 : _GEN_2516; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2518 = 8'hd6 == inBytes_9 ? 8'hf6 : _GEN_2517; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2519 = 8'hd7 == inBytes_9 ? 8'he : _GEN_2518; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2520 = 8'hd8 == inBytes_9 ? 8'h61 : _GEN_2519; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2521 = 8'hd9 == inBytes_9 ? 8'h35 : _GEN_2520; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2522 = 8'hda == inBytes_9 ? 8'h57 : _GEN_2521; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2523 = 8'hdb == inBytes_9 ? 8'hb9 : _GEN_2522; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2524 = 8'hdc == inBytes_9 ? 8'h86 : _GEN_2523; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2525 = 8'hdd == inBytes_9 ? 8'hc1 : _GEN_2524; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2526 = 8'hde == inBytes_9 ? 8'h1d : _GEN_2525; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2527 = 8'hdf == inBytes_9 ? 8'h9e : _GEN_2526; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2528 = 8'he0 == inBytes_9 ? 8'he1 : _GEN_2527; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2529 = 8'he1 == inBytes_9 ? 8'hf8 : _GEN_2528; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2530 = 8'he2 == inBytes_9 ? 8'h98 : _GEN_2529; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2531 = 8'he3 == inBytes_9 ? 8'h11 : _GEN_2530; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2532 = 8'he4 == inBytes_9 ? 8'h69 : _GEN_2531; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2533 = 8'he5 == inBytes_9 ? 8'hd9 : _GEN_2532; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2534 = 8'he6 == inBytes_9 ? 8'h8e : _GEN_2533; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2535 = 8'he7 == inBytes_9 ? 8'h94 : _GEN_2534; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2536 = 8'he8 == inBytes_9 ? 8'h9b : _GEN_2535; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2537 = 8'he9 == inBytes_9 ? 8'h1e : _GEN_2536; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2538 = 8'hea == inBytes_9 ? 8'h87 : _GEN_2537; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2539 = 8'heb == inBytes_9 ? 8'he9 : _GEN_2538; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2540 = 8'hec == inBytes_9 ? 8'hce : _GEN_2539; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2541 = 8'hed == inBytes_9 ? 8'h55 : _GEN_2540; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2542 = 8'hee == inBytes_9 ? 8'h28 : _GEN_2541; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2543 = 8'hef == inBytes_9 ? 8'hdf : _GEN_2542; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2544 = 8'hf0 == inBytes_9 ? 8'h8c : _GEN_2543; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2545 = 8'hf1 == inBytes_9 ? 8'ha1 : _GEN_2544; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2546 = 8'hf2 == inBytes_9 ? 8'h89 : _GEN_2545; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2547 = 8'hf3 == inBytes_9 ? 8'hd : _GEN_2546; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2548 = 8'hf4 == inBytes_9 ? 8'hbf : _GEN_2547; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2549 = 8'hf5 == inBytes_9 ? 8'he6 : _GEN_2548; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2550 = 8'hf6 == inBytes_9 ? 8'h42 : _GEN_2549; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2551 = 8'hf7 == inBytes_9 ? 8'h68 : _GEN_2550; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2552 = 8'hf8 == inBytes_9 ? 8'h41 : _GEN_2551; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2553 = 8'hf9 == inBytes_9 ? 8'h99 : _GEN_2552; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2554 = 8'hfa == inBytes_9 ? 8'h2d : _GEN_2553; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2555 = 8'hfb == inBytes_9 ? 8'hf : _GEN_2554; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2556 = 8'hfc == inBytes_9 ? 8'hb0 : _GEN_2555; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2557 = 8'hfd == inBytes_9 ? 8'h54 : _GEN_2556; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2558 = 8'hfe == inBytes_9 ? 8'hbb : _GEN_2557; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] outBytes_9 = 8'hff == inBytes_9 ? 8'h16 : _GEN_2558; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2561 = 8'h1 == inBytes_10 ? 8'h7c : 8'h63; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2562 = 8'h2 == inBytes_10 ? 8'h77 : _GEN_2561; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2563 = 8'h3 == inBytes_10 ? 8'h7b : _GEN_2562; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2564 = 8'h4 == inBytes_10 ? 8'hf2 : _GEN_2563; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2565 = 8'h5 == inBytes_10 ? 8'h6b : _GEN_2564; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2566 = 8'h6 == inBytes_10 ? 8'h6f : _GEN_2565; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2567 = 8'h7 == inBytes_10 ? 8'hc5 : _GEN_2566; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2568 = 8'h8 == inBytes_10 ? 8'h30 : _GEN_2567; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2569 = 8'h9 == inBytes_10 ? 8'h1 : _GEN_2568; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2570 = 8'ha == inBytes_10 ? 8'h67 : _GEN_2569; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2571 = 8'hb == inBytes_10 ? 8'h2b : _GEN_2570; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2572 = 8'hc == inBytes_10 ? 8'hfe : _GEN_2571; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2573 = 8'hd == inBytes_10 ? 8'hd7 : _GEN_2572; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2574 = 8'he == inBytes_10 ? 8'hab : _GEN_2573; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2575 = 8'hf == inBytes_10 ? 8'h76 : _GEN_2574; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2576 = 8'h10 == inBytes_10 ? 8'hca : _GEN_2575; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2577 = 8'h11 == inBytes_10 ? 8'h82 : _GEN_2576; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2578 = 8'h12 == inBytes_10 ? 8'hc9 : _GEN_2577; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2579 = 8'h13 == inBytes_10 ? 8'h7d : _GEN_2578; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2580 = 8'h14 == inBytes_10 ? 8'hfa : _GEN_2579; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2581 = 8'h15 == inBytes_10 ? 8'h59 : _GEN_2580; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2582 = 8'h16 == inBytes_10 ? 8'h47 : _GEN_2581; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2583 = 8'h17 == inBytes_10 ? 8'hf0 : _GEN_2582; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2584 = 8'h18 == inBytes_10 ? 8'had : _GEN_2583; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2585 = 8'h19 == inBytes_10 ? 8'hd4 : _GEN_2584; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2586 = 8'h1a == inBytes_10 ? 8'ha2 : _GEN_2585; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2587 = 8'h1b == inBytes_10 ? 8'haf : _GEN_2586; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2588 = 8'h1c == inBytes_10 ? 8'h9c : _GEN_2587; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2589 = 8'h1d == inBytes_10 ? 8'ha4 : _GEN_2588; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2590 = 8'h1e == inBytes_10 ? 8'h72 : _GEN_2589; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2591 = 8'h1f == inBytes_10 ? 8'hc0 : _GEN_2590; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2592 = 8'h20 == inBytes_10 ? 8'hb7 : _GEN_2591; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2593 = 8'h21 == inBytes_10 ? 8'hfd : _GEN_2592; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2594 = 8'h22 == inBytes_10 ? 8'h93 : _GEN_2593; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2595 = 8'h23 == inBytes_10 ? 8'h26 : _GEN_2594; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2596 = 8'h24 == inBytes_10 ? 8'h36 : _GEN_2595; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2597 = 8'h25 == inBytes_10 ? 8'h3f : _GEN_2596; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2598 = 8'h26 == inBytes_10 ? 8'hf7 : _GEN_2597; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2599 = 8'h27 == inBytes_10 ? 8'hcc : _GEN_2598; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2600 = 8'h28 == inBytes_10 ? 8'h34 : _GEN_2599; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2601 = 8'h29 == inBytes_10 ? 8'ha5 : _GEN_2600; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2602 = 8'h2a == inBytes_10 ? 8'he5 : _GEN_2601; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2603 = 8'h2b == inBytes_10 ? 8'hf1 : _GEN_2602; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2604 = 8'h2c == inBytes_10 ? 8'h71 : _GEN_2603; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2605 = 8'h2d == inBytes_10 ? 8'hd8 : _GEN_2604; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2606 = 8'h2e == inBytes_10 ? 8'h31 : _GEN_2605; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2607 = 8'h2f == inBytes_10 ? 8'h15 : _GEN_2606; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2608 = 8'h30 == inBytes_10 ? 8'h4 : _GEN_2607; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2609 = 8'h31 == inBytes_10 ? 8'hc7 : _GEN_2608; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2610 = 8'h32 == inBytes_10 ? 8'h23 : _GEN_2609; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2611 = 8'h33 == inBytes_10 ? 8'hc3 : _GEN_2610; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2612 = 8'h34 == inBytes_10 ? 8'h18 : _GEN_2611; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2613 = 8'h35 == inBytes_10 ? 8'h96 : _GEN_2612; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2614 = 8'h36 == inBytes_10 ? 8'h5 : _GEN_2613; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2615 = 8'h37 == inBytes_10 ? 8'h9a : _GEN_2614; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2616 = 8'h38 == inBytes_10 ? 8'h7 : _GEN_2615; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2617 = 8'h39 == inBytes_10 ? 8'h12 : _GEN_2616; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2618 = 8'h3a == inBytes_10 ? 8'h80 : _GEN_2617; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2619 = 8'h3b == inBytes_10 ? 8'he2 : _GEN_2618; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2620 = 8'h3c == inBytes_10 ? 8'heb : _GEN_2619; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2621 = 8'h3d == inBytes_10 ? 8'h27 : _GEN_2620; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2622 = 8'h3e == inBytes_10 ? 8'hb2 : _GEN_2621; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2623 = 8'h3f == inBytes_10 ? 8'h75 : _GEN_2622; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2624 = 8'h40 == inBytes_10 ? 8'h9 : _GEN_2623; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2625 = 8'h41 == inBytes_10 ? 8'h83 : _GEN_2624; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2626 = 8'h42 == inBytes_10 ? 8'h2c : _GEN_2625; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2627 = 8'h43 == inBytes_10 ? 8'h1a : _GEN_2626; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2628 = 8'h44 == inBytes_10 ? 8'h1b : _GEN_2627; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2629 = 8'h45 == inBytes_10 ? 8'h6e : _GEN_2628; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2630 = 8'h46 == inBytes_10 ? 8'h5a : _GEN_2629; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2631 = 8'h47 == inBytes_10 ? 8'ha0 : _GEN_2630; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2632 = 8'h48 == inBytes_10 ? 8'h52 : _GEN_2631; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2633 = 8'h49 == inBytes_10 ? 8'h3b : _GEN_2632; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2634 = 8'h4a == inBytes_10 ? 8'hd6 : _GEN_2633; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2635 = 8'h4b == inBytes_10 ? 8'hb3 : _GEN_2634; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2636 = 8'h4c == inBytes_10 ? 8'h29 : _GEN_2635; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2637 = 8'h4d == inBytes_10 ? 8'he3 : _GEN_2636; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2638 = 8'h4e == inBytes_10 ? 8'h2f : _GEN_2637; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2639 = 8'h4f == inBytes_10 ? 8'h84 : _GEN_2638; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2640 = 8'h50 == inBytes_10 ? 8'h53 : _GEN_2639; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2641 = 8'h51 == inBytes_10 ? 8'hd1 : _GEN_2640; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2642 = 8'h52 == inBytes_10 ? 8'h0 : _GEN_2641; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2643 = 8'h53 == inBytes_10 ? 8'hed : _GEN_2642; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2644 = 8'h54 == inBytes_10 ? 8'h20 : _GEN_2643; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2645 = 8'h55 == inBytes_10 ? 8'hfc : _GEN_2644; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2646 = 8'h56 == inBytes_10 ? 8'hb1 : _GEN_2645; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2647 = 8'h57 == inBytes_10 ? 8'h5b : _GEN_2646; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2648 = 8'h58 == inBytes_10 ? 8'h6a : _GEN_2647; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2649 = 8'h59 == inBytes_10 ? 8'hcb : _GEN_2648; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2650 = 8'h5a == inBytes_10 ? 8'hbe : _GEN_2649; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2651 = 8'h5b == inBytes_10 ? 8'h39 : _GEN_2650; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2652 = 8'h5c == inBytes_10 ? 8'h4a : _GEN_2651; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2653 = 8'h5d == inBytes_10 ? 8'h4c : _GEN_2652; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2654 = 8'h5e == inBytes_10 ? 8'h58 : _GEN_2653; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2655 = 8'h5f == inBytes_10 ? 8'hcf : _GEN_2654; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2656 = 8'h60 == inBytes_10 ? 8'hd0 : _GEN_2655; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2657 = 8'h61 == inBytes_10 ? 8'hef : _GEN_2656; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2658 = 8'h62 == inBytes_10 ? 8'haa : _GEN_2657; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2659 = 8'h63 == inBytes_10 ? 8'hfb : _GEN_2658; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2660 = 8'h64 == inBytes_10 ? 8'h43 : _GEN_2659; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2661 = 8'h65 == inBytes_10 ? 8'h4d : _GEN_2660; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2662 = 8'h66 == inBytes_10 ? 8'h33 : _GEN_2661; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2663 = 8'h67 == inBytes_10 ? 8'h85 : _GEN_2662; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2664 = 8'h68 == inBytes_10 ? 8'h45 : _GEN_2663; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2665 = 8'h69 == inBytes_10 ? 8'hf9 : _GEN_2664; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2666 = 8'h6a == inBytes_10 ? 8'h2 : _GEN_2665; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2667 = 8'h6b == inBytes_10 ? 8'h7f : _GEN_2666; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2668 = 8'h6c == inBytes_10 ? 8'h50 : _GEN_2667; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2669 = 8'h6d == inBytes_10 ? 8'h3c : _GEN_2668; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2670 = 8'h6e == inBytes_10 ? 8'h9f : _GEN_2669; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2671 = 8'h6f == inBytes_10 ? 8'ha8 : _GEN_2670; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2672 = 8'h70 == inBytes_10 ? 8'h51 : _GEN_2671; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2673 = 8'h71 == inBytes_10 ? 8'ha3 : _GEN_2672; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2674 = 8'h72 == inBytes_10 ? 8'h40 : _GEN_2673; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2675 = 8'h73 == inBytes_10 ? 8'h8f : _GEN_2674; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2676 = 8'h74 == inBytes_10 ? 8'h92 : _GEN_2675; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2677 = 8'h75 == inBytes_10 ? 8'h9d : _GEN_2676; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2678 = 8'h76 == inBytes_10 ? 8'h38 : _GEN_2677; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2679 = 8'h77 == inBytes_10 ? 8'hf5 : _GEN_2678; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2680 = 8'h78 == inBytes_10 ? 8'hbc : _GEN_2679; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2681 = 8'h79 == inBytes_10 ? 8'hb6 : _GEN_2680; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2682 = 8'h7a == inBytes_10 ? 8'hda : _GEN_2681; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2683 = 8'h7b == inBytes_10 ? 8'h21 : _GEN_2682; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2684 = 8'h7c == inBytes_10 ? 8'h10 : _GEN_2683; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2685 = 8'h7d == inBytes_10 ? 8'hff : _GEN_2684; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2686 = 8'h7e == inBytes_10 ? 8'hf3 : _GEN_2685; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2687 = 8'h7f == inBytes_10 ? 8'hd2 : _GEN_2686; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2688 = 8'h80 == inBytes_10 ? 8'hcd : _GEN_2687; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2689 = 8'h81 == inBytes_10 ? 8'hc : _GEN_2688; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2690 = 8'h82 == inBytes_10 ? 8'h13 : _GEN_2689; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2691 = 8'h83 == inBytes_10 ? 8'hec : _GEN_2690; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2692 = 8'h84 == inBytes_10 ? 8'h5f : _GEN_2691; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2693 = 8'h85 == inBytes_10 ? 8'h97 : _GEN_2692; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2694 = 8'h86 == inBytes_10 ? 8'h44 : _GEN_2693; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2695 = 8'h87 == inBytes_10 ? 8'h17 : _GEN_2694; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2696 = 8'h88 == inBytes_10 ? 8'hc4 : _GEN_2695; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2697 = 8'h89 == inBytes_10 ? 8'ha7 : _GEN_2696; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2698 = 8'h8a == inBytes_10 ? 8'h7e : _GEN_2697; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2699 = 8'h8b == inBytes_10 ? 8'h3d : _GEN_2698; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2700 = 8'h8c == inBytes_10 ? 8'h64 : _GEN_2699; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2701 = 8'h8d == inBytes_10 ? 8'h5d : _GEN_2700; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2702 = 8'h8e == inBytes_10 ? 8'h19 : _GEN_2701; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2703 = 8'h8f == inBytes_10 ? 8'h73 : _GEN_2702; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2704 = 8'h90 == inBytes_10 ? 8'h60 : _GEN_2703; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2705 = 8'h91 == inBytes_10 ? 8'h81 : _GEN_2704; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2706 = 8'h92 == inBytes_10 ? 8'h4f : _GEN_2705; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2707 = 8'h93 == inBytes_10 ? 8'hdc : _GEN_2706; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2708 = 8'h94 == inBytes_10 ? 8'h22 : _GEN_2707; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2709 = 8'h95 == inBytes_10 ? 8'h2a : _GEN_2708; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2710 = 8'h96 == inBytes_10 ? 8'h90 : _GEN_2709; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2711 = 8'h97 == inBytes_10 ? 8'h88 : _GEN_2710; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2712 = 8'h98 == inBytes_10 ? 8'h46 : _GEN_2711; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2713 = 8'h99 == inBytes_10 ? 8'hee : _GEN_2712; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2714 = 8'h9a == inBytes_10 ? 8'hb8 : _GEN_2713; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2715 = 8'h9b == inBytes_10 ? 8'h14 : _GEN_2714; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2716 = 8'h9c == inBytes_10 ? 8'hde : _GEN_2715; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2717 = 8'h9d == inBytes_10 ? 8'h5e : _GEN_2716; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2718 = 8'h9e == inBytes_10 ? 8'hb : _GEN_2717; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2719 = 8'h9f == inBytes_10 ? 8'hdb : _GEN_2718; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2720 = 8'ha0 == inBytes_10 ? 8'he0 : _GEN_2719; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2721 = 8'ha1 == inBytes_10 ? 8'h32 : _GEN_2720; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2722 = 8'ha2 == inBytes_10 ? 8'h3a : _GEN_2721; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2723 = 8'ha3 == inBytes_10 ? 8'ha : _GEN_2722; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2724 = 8'ha4 == inBytes_10 ? 8'h49 : _GEN_2723; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2725 = 8'ha5 == inBytes_10 ? 8'h6 : _GEN_2724; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2726 = 8'ha6 == inBytes_10 ? 8'h24 : _GEN_2725; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2727 = 8'ha7 == inBytes_10 ? 8'h5c : _GEN_2726; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2728 = 8'ha8 == inBytes_10 ? 8'hc2 : _GEN_2727; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2729 = 8'ha9 == inBytes_10 ? 8'hd3 : _GEN_2728; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2730 = 8'haa == inBytes_10 ? 8'hac : _GEN_2729; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2731 = 8'hab == inBytes_10 ? 8'h62 : _GEN_2730; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2732 = 8'hac == inBytes_10 ? 8'h91 : _GEN_2731; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2733 = 8'had == inBytes_10 ? 8'h95 : _GEN_2732; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2734 = 8'hae == inBytes_10 ? 8'he4 : _GEN_2733; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2735 = 8'haf == inBytes_10 ? 8'h79 : _GEN_2734; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2736 = 8'hb0 == inBytes_10 ? 8'he7 : _GEN_2735; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2737 = 8'hb1 == inBytes_10 ? 8'hc8 : _GEN_2736; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2738 = 8'hb2 == inBytes_10 ? 8'h37 : _GEN_2737; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2739 = 8'hb3 == inBytes_10 ? 8'h6d : _GEN_2738; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2740 = 8'hb4 == inBytes_10 ? 8'h8d : _GEN_2739; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2741 = 8'hb5 == inBytes_10 ? 8'hd5 : _GEN_2740; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2742 = 8'hb6 == inBytes_10 ? 8'h4e : _GEN_2741; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2743 = 8'hb7 == inBytes_10 ? 8'ha9 : _GEN_2742; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2744 = 8'hb8 == inBytes_10 ? 8'h6c : _GEN_2743; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2745 = 8'hb9 == inBytes_10 ? 8'h56 : _GEN_2744; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2746 = 8'hba == inBytes_10 ? 8'hf4 : _GEN_2745; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2747 = 8'hbb == inBytes_10 ? 8'hea : _GEN_2746; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2748 = 8'hbc == inBytes_10 ? 8'h65 : _GEN_2747; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2749 = 8'hbd == inBytes_10 ? 8'h7a : _GEN_2748; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2750 = 8'hbe == inBytes_10 ? 8'hae : _GEN_2749; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2751 = 8'hbf == inBytes_10 ? 8'h8 : _GEN_2750; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2752 = 8'hc0 == inBytes_10 ? 8'hba : _GEN_2751; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2753 = 8'hc1 == inBytes_10 ? 8'h78 : _GEN_2752; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2754 = 8'hc2 == inBytes_10 ? 8'h25 : _GEN_2753; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2755 = 8'hc3 == inBytes_10 ? 8'h2e : _GEN_2754; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2756 = 8'hc4 == inBytes_10 ? 8'h1c : _GEN_2755; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2757 = 8'hc5 == inBytes_10 ? 8'ha6 : _GEN_2756; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2758 = 8'hc6 == inBytes_10 ? 8'hb4 : _GEN_2757; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2759 = 8'hc7 == inBytes_10 ? 8'hc6 : _GEN_2758; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2760 = 8'hc8 == inBytes_10 ? 8'he8 : _GEN_2759; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2761 = 8'hc9 == inBytes_10 ? 8'hdd : _GEN_2760; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2762 = 8'hca == inBytes_10 ? 8'h74 : _GEN_2761; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2763 = 8'hcb == inBytes_10 ? 8'h1f : _GEN_2762; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2764 = 8'hcc == inBytes_10 ? 8'h4b : _GEN_2763; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2765 = 8'hcd == inBytes_10 ? 8'hbd : _GEN_2764; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2766 = 8'hce == inBytes_10 ? 8'h8b : _GEN_2765; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2767 = 8'hcf == inBytes_10 ? 8'h8a : _GEN_2766; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2768 = 8'hd0 == inBytes_10 ? 8'h70 : _GEN_2767; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2769 = 8'hd1 == inBytes_10 ? 8'h3e : _GEN_2768; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2770 = 8'hd2 == inBytes_10 ? 8'hb5 : _GEN_2769; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2771 = 8'hd3 == inBytes_10 ? 8'h66 : _GEN_2770; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2772 = 8'hd4 == inBytes_10 ? 8'h48 : _GEN_2771; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2773 = 8'hd5 == inBytes_10 ? 8'h3 : _GEN_2772; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2774 = 8'hd6 == inBytes_10 ? 8'hf6 : _GEN_2773; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2775 = 8'hd7 == inBytes_10 ? 8'he : _GEN_2774; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2776 = 8'hd8 == inBytes_10 ? 8'h61 : _GEN_2775; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2777 = 8'hd9 == inBytes_10 ? 8'h35 : _GEN_2776; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2778 = 8'hda == inBytes_10 ? 8'h57 : _GEN_2777; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2779 = 8'hdb == inBytes_10 ? 8'hb9 : _GEN_2778; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2780 = 8'hdc == inBytes_10 ? 8'h86 : _GEN_2779; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2781 = 8'hdd == inBytes_10 ? 8'hc1 : _GEN_2780; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2782 = 8'hde == inBytes_10 ? 8'h1d : _GEN_2781; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2783 = 8'hdf == inBytes_10 ? 8'h9e : _GEN_2782; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2784 = 8'he0 == inBytes_10 ? 8'he1 : _GEN_2783; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2785 = 8'he1 == inBytes_10 ? 8'hf8 : _GEN_2784; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2786 = 8'he2 == inBytes_10 ? 8'h98 : _GEN_2785; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2787 = 8'he3 == inBytes_10 ? 8'h11 : _GEN_2786; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2788 = 8'he4 == inBytes_10 ? 8'h69 : _GEN_2787; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2789 = 8'he5 == inBytes_10 ? 8'hd9 : _GEN_2788; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2790 = 8'he6 == inBytes_10 ? 8'h8e : _GEN_2789; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2791 = 8'he7 == inBytes_10 ? 8'h94 : _GEN_2790; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2792 = 8'he8 == inBytes_10 ? 8'h9b : _GEN_2791; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2793 = 8'he9 == inBytes_10 ? 8'h1e : _GEN_2792; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2794 = 8'hea == inBytes_10 ? 8'h87 : _GEN_2793; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2795 = 8'heb == inBytes_10 ? 8'he9 : _GEN_2794; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2796 = 8'hec == inBytes_10 ? 8'hce : _GEN_2795; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2797 = 8'hed == inBytes_10 ? 8'h55 : _GEN_2796; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2798 = 8'hee == inBytes_10 ? 8'h28 : _GEN_2797; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2799 = 8'hef == inBytes_10 ? 8'hdf : _GEN_2798; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2800 = 8'hf0 == inBytes_10 ? 8'h8c : _GEN_2799; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2801 = 8'hf1 == inBytes_10 ? 8'ha1 : _GEN_2800; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2802 = 8'hf2 == inBytes_10 ? 8'h89 : _GEN_2801; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2803 = 8'hf3 == inBytes_10 ? 8'hd : _GEN_2802; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2804 = 8'hf4 == inBytes_10 ? 8'hbf : _GEN_2803; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2805 = 8'hf5 == inBytes_10 ? 8'he6 : _GEN_2804; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2806 = 8'hf6 == inBytes_10 ? 8'h42 : _GEN_2805; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2807 = 8'hf7 == inBytes_10 ? 8'h68 : _GEN_2806; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2808 = 8'hf8 == inBytes_10 ? 8'h41 : _GEN_2807; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2809 = 8'hf9 == inBytes_10 ? 8'h99 : _GEN_2808; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2810 = 8'hfa == inBytes_10 ? 8'h2d : _GEN_2809; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2811 = 8'hfb == inBytes_10 ? 8'hf : _GEN_2810; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2812 = 8'hfc == inBytes_10 ? 8'hb0 : _GEN_2811; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2813 = 8'hfd == inBytes_10 ? 8'h54 : _GEN_2812; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2814 = 8'hfe == inBytes_10 ? 8'hbb : _GEN_2813; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] outBytes_10 = 8'hff == inBytes_10 ? 8'h16 : _GEN_2814; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2817 = 8'h1 == inBytes_11 ? 8'h7c : 8'h63; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2818 = 8'h2 == inBytes_11 ? 8'h77 : _GEN_2817; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2819 = 8'h3 == inBytes_11 ? 8'h7b : _GEN_2818; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2820 = 8'h4 == inBytes_11 ? 8'hf2 : _GEN_2819; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2821 = 8'h5 == inBytes_11 ? 8'h6b : _GEN_2820; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2822 = 8'h6 == inBytes_11 ? 8'h6f : _GEN_2821; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2823 = 8'h7 == inBytes_11 ? 8'hc5 : _GEN_2822; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2824 = 8'h8 == inBytes_11 ? 8'h30 : _GEN_2823; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2825 = 8'h9 == inBytes_11 ? 8'h1 : _GEN_2824; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2826 = 8'ha == inBytes_11 ? 8'h67 : _GEN_2825; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2827 = 8'hb == inBytes_11 ? 8'h2b : _GEN_2826; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2828 = 8'hc == inBytes_11 ? 8'hfe : _GEN_2827; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2829 = 8'hd == inBytes_11 ? 8'hd7 : _GEN_2828; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2830 = 8'he == inBytes_11 ? 8'hab : _GEN_2829; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2831 = 8'hf == inBytes_11 ? 8'h76 : _GEN_2830; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2832 = 8'h10 == inBytes_11 ? 8'hca : _GEN_2831; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2833 = 8'h11 == inBytes_11 ? 8'h82 : _GEN_2832; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2834 = 8'h12 == inBytes_11 ? 8'hc9 : _GEN_2833; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2835 = 8'h13 == inBytes_11 ? 8'h7d : _GEN_2834; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2836 = 8'h14 == inBytes_11 ? 8'hfa : _GEN_2835; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2837 = 8'h15 == inBytes_11 ? 8'h59 : _GEN_2836; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2838 = 8'h16 == inBytes_11 ? 8'h47 : _GEN_2837; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2839 = 8'h17 == inBytes_11 ? 8'hf0 : _GEN_2838; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2840 = 8'h18 == inBytes_11 ? 8'had : _GEN_2839; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2841 = 8'h19 == inBytes_11 ? 8'hd4 : _GEN_2840; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2842 = 8'h1a == inBytes_11 ? 8'ha2 : _GEN_2841; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2843 = 8'h1b == inBytes_11 ? 8'haf : _GEN_2842; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2844 = 8'h1c == inBytes_11 ? 8'h9c : _GEN_2843; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2845 = 8'h1d == inBytes_11 ? 8'ha4 : _GEN_2844; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2846 = 8'h1e == inBytes_11 ? 8'h72 : _GEN_2845; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2847 = 8'h1f == inBytes_11 ? 8'hc0 : _GEN_2846; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2848 = 8'h20 == inBytes_11 ? 8'hb7 : _GEN_2847; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2849 = 8'h21 == inBytes_11 ? 8'hfd : _GEN_2848; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2850 = 8'h22 == inBytes_11 ? 8'h93 : _GEN_2849; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2851 = 8'h23 == inBytes_11 ? 8'h26 : _GEN_2850; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2852 = 8'h24 == inBytes_11 ? 8'h36 : _GEN_2851; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2853 = 8'h25 == inBytes_11 ? 8'h3f : _GEN_2852; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2854 = 8'h26 == inBytes_11 ? 8'hf7 : _GEN_2853; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2855 = 8'h27 == inBytes_11 ? 8'hcc : _GEN_2854; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2856 = 8'h28 == inBytes_11 ? 8'h34 : _GEN_2855; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2857 = 8'h29 == inBytes_11 ? 8'ha5 : _GEN_2856; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2858 = 8'h2a == inBytes_11 ? 8'he5 : _GEN_2857; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2859 = 8'h2b == inBytes_11 ? 8'hf1 : _GEN_2858; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2860 = 8'h2c == inBytes_11 ? 8'h71 : _GEN_2859; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2861 = 8'h2d == inBytes_11 ? 8'hd8 : _GEN_2860; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2862 = 8'h2e == inBytes_11 ? 8'h31 : _GEN_2861; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2863 = 8'h2f == inBytes_11 ? 8'h15 : _GEN_2862; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2864 = 8'h30 == inBytes_11 ? 8'h4 : _GEN_2863; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2865 = 8'h31 == inBytes_11 ? 8'hc7 : _GEN_2864; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2866 = 8'h32 == inBytes_11 ? 8'h23 : _GEN_2865; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2867 = 8'h33 == inBytes_11 ? 8'hc3 : _GEN_2866; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2868 = 8'h34 == inBytes_11 ? 8'h18 : _GEN_2867; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2869 = 8'h35 == inBytes_11 ? 8'h96 : _GEN_2868; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2870 = 8'h36 == inBytes_11 ? 8'h5 : _GEN_2869; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2871 = 8'h37 == inBytes_11 ? 8'h9a : _GEN_2870; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2872 = 8'h38 == inBytes_11 ? 8'h7 : _GEN_2871; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2873 = 8'h39 == inBytes_11 ? 8'h12 : _GEN_2872; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2874 = 8'h3a == inBytes_11 ? 8'h80 : _GEN_2873; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2875 = 8'h3b == inBytes_11 ? 8'he2 : _GEN_2874; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2876 = 8'h3c == inBytes_11 ? 8'heb : _GEN_2875; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2877 = 8'h3d == inBytes_11 ? 8'h27 : _GEN_2876; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2878 = 8'h3e == inBytes_11 ? 8'hb2 : _GEN_2877; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2879 = 8'h3f == inBytes_11 ? 8'h75 : _GEN_2878; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2880 = 8'h40 == inBytes_11 ? 8'h9 : _GEN_2879; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2881 = 8'h41 == inBytes_11 ? 8'h83 : _GEN_2880; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2882 = 8'h42 == inBytes_11 ? 8'h2c : _GEN_2881; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2883 = 8'h43 == inBytes_11 ? 8'h1a : _GEN_2882; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2884 = 8'h44 == inBytes_11 ? 8'h1b : _GEN_2883; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2885 = 8'h45 == inBytes_11 ? 8'h6e : _GEN_2884; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2886 = 8'h46 == inBytes_11 ? 8'h5a : _GEN_2885; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2887 = 8'h47 == inBytes_11 ? 8'ha0 : _GEN_2886; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2888 = 8'h48 == inBytes_11 ? 8'h52 : _GEN_2887; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2889 = 8'h49 == inBytes_11 ? 8'h3b : _GEN_2888; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2890 = 8'h4a == inBytes_11 ? 8'hd6 : _GEN_2889; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2891 = 8'h4b == inBytes_11 ? 8'hb3 : _GEN_2890; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2892 = 8'h4c == inBytes_11 ? 8'h29 : _GEN_2891; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2893 = 8'h4d == inBytes_11 ? 8'he3 : _GEN_2892; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2894 = 8'h4e == inBytes_11 ? 8'h2f : _GEN_2893; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2895 = 8'h4f == inBytes_11 ? 8'h84 : _GEN_2894; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2896 = 8'h50 == inBytes_11 ? 8'h53 : _GEN_2895; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2897 = 8'h51 == inBytes_11 ? 8'hd1 : _GEN_2896; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2898 = 8'h52 == inBytes_11 ? 8'h0 : _GEN_2897; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2899 = 8'h53 == inBytes_11 ? 8'hed : _GEN_2898; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2900 = 8'h54 == inBytes_11 ? 8'h20 : _GEN_2899; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2901 = 8'h55 == inBytes_11 ? 8'hfc : _GEN_2900; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2902 = 8'h56 == inBytes_11 ? 8'hb1 : _GEN_2901; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2903 = 8'h57 == inBytes_11 ? 8'h5b : _GEN_2902; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2904 = 8'h58 == inBytes_11 ? 8'h6a : _GEN_2903; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2905 = 8'h59 == inBytes_11 ? 8'hcb : _GEN_2904; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2906 = 8'h5a == inBytes_11 ? 8'hbe : _GEN_2905; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2907 = 8'h5b == inBytes_11 ? 8'h39 : _GEN_2906; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2908 = 8'h5c == inBytes_11 ? 8'h4a : _GEN_2907; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2909 = 8'h5d == inBytes_11 ? 8'h4c : _GEN_2908; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2910 = 8'h5e == inBytes_11 ? 8'h58 : _GEN_2909; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2911 = 8'h5f == inBytes_11 ? 8'hcf : _GEN_2910; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2912 = 8'h60 == inBytes_11 ? 8'hd0 : _GEN_2911; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2913 = 8'h61 == inBytes_11 ? 8'hef : _GEN_2912; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2914 = 8'h62 == inBytes_11 ? 8'haa : _GEN_2913; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2915 = 8'h63 == inBytes_11 ? 8'hfb : _GEN_2914; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2916 = 8'h64 == inBytes_11 ? 8'h43 : _GEN_2915; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2917 = 8'h65 == inBytes_11 ? 8'h4d : _GEN_2916; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2918 = 8'h66 == inBytes_11 ? 8'h33 : _GEN_2917; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2919 = 8'h67 == inBytes_11 ? 8'h85 : _GEN_2918; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2920 = 8'h68 == inBytes_11 ? 8'h45 : _GEN_2919; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2921 = 8'h69 == inBytes_11 ? 8'hf9 : _GEN_2920; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2922 = 8'h6a == inBytes_11 ? 8'h2 : _GEN_2921; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2923 = 8'h6b == inBytes_11 ? 8'h7f : _GEN_2922; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2924 = 8'h6c == inBytes_11 ? 8'h50 : _GEN_2923; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2925 = 8'h6d == inBytes_11 ? 8'h3c : _GEN_2924; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2926 = 8'h6e == inBytes_11 ? 8'h9f : _GEN_2925; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2927 = 8'h6f == inBytes_11 ? 8'ha8 : _GEN_2926; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2928 = 8'h70 == inBytes_11 ? 8'h51 : _GEN_2927; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2929 = 8'h71 == inBytes_11 ? 8'ha3 : _GEN_2928; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2930 = 8'h72 == inBytes_11 ? 8'h40 : _GEN_2929; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2931 = 8'h73 == inBytes_11 ? 8'h8f : _GEN_2930; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2932 = 8'h74 == inBytes_11 ? 8'h92 : _GEN_2931; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2933 = 8'h75 == inBytes_11 ? 8'h9d : _GEN_2932; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2934 = 8'h76 == inBytes_11 ? 8'h38 : _GEN_2933; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2935 = 8'h77 == inBytes_11 ? 8'hf5 : _GEN_2934; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2936 = 8'h78 == inBytes_11 ? 8'hbc : _GEN_2935; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2937 = 8'h79 == inBytes_11 ? 8'hb6 : _GEN_2936; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2938 = 8'h7a == inBytes_11 ? 8'hda : _GEN_2937; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2939 = 8'h7b == inBytes_11 ? 8'h21 : _GEN_2938; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2940 = 8'h7c == inBytes_11 ? 8'h10 : _GEN_2939; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2941 = 8'h7d == inBytes_11 ? 8'hff : _GEN_2940; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2942 = 8'h7e == inBytes_11 ? 8'hf3 : _GEN_2941; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2943 = 8'h7f == inBytes_11 ? 8'hd2 : _GEN_2942; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2944 = 8'h80 == inBytes_11 ? 8'hcd : _GEN_2943; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2945 = 8'h81 == inBytes_11 ? 8'hc : _GEN_2944; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2946 = 8'h82 == inBytes_11 ? 8'h13 : _GEN_2945; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2947 = 8'h83 == inBytes_11 ? 8'hec : _GEN_2946; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2948 = 8'h84 == inBytes_11 ? 8'h5f : _GEN_2947; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2949 = 8'h85 == inBytes_11 ? 8'h97 : _GEN_2948; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2950 = 8'h86 == inBytes_11 ? 8'h44 : _GEN_2949; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2951 = 8'h87 == inBytes_11 ? 8'h17 : _GEN_2950; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2952 = 8'h88 == inBytes_11 ? 8'hc4 : _GEN_2951; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2953 = 8'h89 == inBytes_11 ? 8'ha7 : _GEN_2952; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2954 = 8'h8a == inBytes_11 ? 8'h7e : _GEN_2953; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2955 = 8'h8b == inBytes_11 ? 8'h3d : _GEN_2954; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2956 = 8'h8c == inBytes_11 ? 8'h64 : _GEN_2955; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2957 = 8'h8d == inBytes_11 ? 8'h5d : _GEN_2956; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2958 = 8'h8e == inBytes_11 ? 8'h19 : _GEN_2957; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2959 = 8'h8f == inBytes_11 ? 8'h73 : _GEN_2958; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2960 = 8'h90 == inBytes_11 ? 8'h60 : _GEN_2959; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2961 = 8'h91 == inBytes_11 ? 8'h81 : _GEN_2960; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2962 = 8'h92 == inBytes_11 ? 8'h4f : _GEN_2961; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2963 = 8'h93 == inBytes_11 ? 8'hdc : _GEN_2962; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2964 = 8'h94 == inBytes_11 ? 8'h22 : _GEN_2963; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2965 = 8'h95 == inBytes_11 ? 8'h2a : _GEN_2964; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2966 = 8'h96 == inBytes_11 ? 8'h90 : _GEN_2965; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2967 = 8'h97 == inBytes_11 ? 8'h88 : _GEN_2966; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2968 = 8'h98 == inBytes_11 ? 8'h46 : _GEN_2967; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2969 = 8'h99 == inBytes_11 ? 8'hee : _GEN_2968; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2970 = 8'h9a == inBytes_11 ? 8'hb8 : _GEN_2969; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2971 = 8'h9b == inBytes_11 ? 8'h14 : _GEN_2970; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2972 = 8'h9c == inBytes_11 ? 8'hde : _GEN_2971; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2973 = 8'h9d == inBytes_11 ? 8'h5e : _GEN_2972; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2974 = 8'h9e == inBytes_11 ? 8'hb : _GEN_2973; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2975 = 8'h9f == inBytes_11 ? 8'hdb : _GEN_2974; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2976 = 8'ha0 == inBytes_11 ? 8'he0 : _GEN_2975; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2977 = 8'ha1 == inBytes_11 ? 8'h32 : _GEN_2976; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2978 = 8'ha2 == inBytes_11 ? 8'h3a : _GEN_2977; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2979 = 8'ha3 == inBytes_11 ? 8'ha : _GEN_2978; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2980 = 8'ha4 == inBytes_11 ? 8'h49 : _GEN_2979; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2981 = 8'ha5 == inBytes_11 ? 8'h6 : _GEN_2980; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2982 = 8'ha6 == inBytes_11 ? 8'h24 : _GEN_2981; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2983 = 8'ha7 == inBytes_11 ? 8'h5c : _GEN_2982; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2984 = 8'ha8 == inBytes_11 ? 8'hc2 : _GEN_2983; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2985 = 8'ha9 == inBytes_11 ? 8'hd3 : _GEN_2984; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2986 = 8'haa == inBytes_11 ? 8'hac : _GEN_2985; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2987 = 8'hab == inBytes_11 ? 8'h62 : _GEN_2986; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2988 = 8'hac == inBytes_11 ? 8'h91 : _GEN_2987; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2989 = 8'had == inBytes_11 ? 8'h95 : _GEN_2988; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2990 = 8'hae == inBytes_11 ? 8'he4 : _GEN_2989; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2991 = 8'haf == inBytes_11 ? 8'h79 : _GEN_2990; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2992 = 8'hb0 == inBytes_11 ? 8'he7 : _GEN_2991; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2993 = 8'hb1 == inBytes_11 ? 8'hc8 : _GEN_2992; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2994 = 8'hb2 == inBytes_11 ? 8'h37 : _GEN_2993; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2995 = 8'hb3 == inBytes_11 ? 8'h6d : _GEN_2994; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2996 = 8'hb4 == inBytes_11 ? 8'h8d : _GEN_2995; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2997 = 8'hb5 == inBytes_11 ? 8'hd5 : _GEN_2996; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2998 = 8'hb6 == inBytes_11 ? 8'h4e : _GEN_2997; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_2999 = 8'hb7 == inBytes_11 ? 8'ha9 : _GEN_2998; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3000 = 8'hb8 == inBytes_11 ? 8'h6c : _GEN_2999; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3001 = 8'hb9 == inBytes_11 ? 8'h56 : _GEN_3000; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3002 = 8'hba == inBytes_11 ? 8'hf4 : _GEN_3001; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3003 = 8'hbb == inBytes_11 ? 8'hea : _GEN_3002; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3004 = 8'hbc == inBytes_11 ? 8'h65 : _GEN_3003; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3005 = 8'hbd == inBytes_11 ? 8'h7a : _GEN_3004; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3006 = 8'hbe == inBytes_11 ? 8'hae : _GEN_3005; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3007 = 8'hbf == inBytes_11 ? 8'h8 : _GEN_3006; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3008 = 8'hc0 == inBytes_11 ? 8'hba : _GEN_3007; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3009 = 8'hc1 == inBytes_11 ? 8'h78 : _GEN_3008; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3010 = 8'hc2 == inBytes_11 ? 8'h25 : _GEN_3009; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3011 = 8'hc3 == inBytes_11 ? 8'h2e : _GEN_3010; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3012 = 8'hc4 == inBytes_11 ? 8'h1c : _GEN_3011; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3013 = 8'hc5 == inBytes_11 ? 8'ha6 : _GEN_3012; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3014 = 8'hc6 == inBytes_11 ? 8'hb4 : _GEN_3013; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3015 = 8'hc7 == inBytes_11 ? 8'hc6 : _GEN_3014; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3016 = 8'hc8 == inBytes_11 ? 8'he8 : _GEN_3015; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3017 = 8'hc9 == inBytes_11 ? 8'hdd : _GEN_3016; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3018 = 8'hca == inBytes_11 ? 8'h74 : _GEN_3017; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3019 = 8'hcb == inBytes_11 ? 8'h1f : _GEN_3018; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3020 = 8'hcc == inBytes_11 ? 8'h4b : _GEN_3019; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3021 = 8'hcd == inBytes_11 ? 8'hbd : _GEN_3020; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3022 = 8'hce == inBytes_11 ? 8'h8b : _GEN_3021; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3023 = 8'hcf == inBytes_11 ? 8'h8a : _GEN_3022; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3024 = 8'hd0 == inBytes_11 ? 8'h70 : _GEN_3023; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3025 = 8'hd1 == inBytes_11 ? 8'h3e : _GEN_3024; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3026 = 8'hd2 == inBytes_11 ? 8'hb5 : _GEN_3025; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3027 = 8'hd3 == inBytes_11 ? 8'h66 : _GEN_3026; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3028 = 8'hd4 == inBytes_11 ? 8'h48 : _GEN_3027; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3029 = 8'hd5 == inBytes_11 ? 8'h3 : _GEN_3028; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3030 = 8'hd6 == inBytes_11 ? 8'hf6 : _GEN_3029; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3031 = 8'hd7 == inBytes_11 ? 8'he : _GEN_3030; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3032 = 8'hd8 == inBytes_11 ? 8'h61 : _GEN_3031; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3033 = 8'hd9 == inBytes_11 ? 8'h35 : _GEN_3032; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3034 = 8'hda == inBytes_11 ? 8'h57 : _GEN_3033; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3035 = 8'hdb == inBytes_11 ? 8'hb9 : _GEN_3034; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3036 = 8'hdc == inBytes_11 ? 8'h86 : _GEN_3035; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3037 = 8'hdd == inBytes_11 ? 8'hc1 : _GEN_3036; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3038 = 8'hde == inBytes_11 ? 8'h1d : _GEN_3037; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3039 = 8'hdf == inBytes_11 ? 8'h9e : _GEN_3038; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3040 = 8'he0 == inBytes_11 ? 8'he1 : _GEN_3039; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3041 = 8'he1 == inBytes_11 ? 8'hf8 : _GEN_3040; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3042 = 8'he2 == inBytes_11 ? 8'h98 : _GEN_3041; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3043 = 8'he3 == inBytes_11 ? 8'h11 : _GEN_3042; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3044 = 8'he4 == inBytes_11 ? 8'h69 : _GEN_3043; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3045 = 8'he5 == inBytes_11 ? 8'hd9 : _GEN_3044; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3046 = 8'he6 == inBytes_11 ? 8'h8e : _GEN_3045; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3047 = 8'he7 == inBytes_11 ? 8'h94 : _GEN_3046; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3048 = 8'he8 == inBytes_11 ? 8'h9b : _GEN_3047; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3049 = 8'he9 == inBytes_11 ? 8'h1e : _GEN_3048; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3050 = 8'hea == inBytes_11 ? 8'h87 : _GEN_3049; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3051 = 8'heb == inBytes_11 ? 8'he9 : _GEN_3050; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3052 = 8'hec == inBytes_11 ? 8'hce : _GEN_3051; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3053 = 8'hed == inBytes_11 ? 8'h55 : _GEN_3052; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3054 = 8'hee == inBytes_11 ? 8'h28 : _GEN_3053; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3055 = 8'hef == inBytes_11 ? 8'hdf : _GEN_3054; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3056 = 8'hf0 == inBytes_11 ? 8'h8c : _GEN_3055; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3057 = 8'hf1 == inBytes_11 ? 8'ha1 : _GEN_3056; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3058 = 8'hf2 == inBytes_11 ? 8'h89 : _GEN_3057; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3059 = 8'hf3 == inBytes_11 ? 8'hd : _GEN_3058; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3060 = 8'hf4 == inBytes_11 ? 8'hbf : _GEN_3059; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3061 = 8'hf5 == inBytes_11 ? 8'he6 : _GEN_3060; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3062 = 8'hf6 == inBytes_11 ? 8'h42 : _GEN_3061; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3063 = 8'hf7 == inBytes_11 ? 8'h68 : _GEN_3062; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3064 = 8'hf8 == inBytes_11 ? 8'h41 : _GEN_3063; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3065 = 8'hf9 == inBytes_11 ? 8'h99 : _GEN_3064; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3066 = 8'hfa == inBytes_11 ? 8'h2d : _GEN_3065; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3067 = 8'hfb == inBytes_11 ? 8'hf : _GEN_3066; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3068 = 8'hfc == inBytes_11 ? 8'hb0 : _GEN_3067; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3069 = 8'hfd == inBytes_11 ? 8'h54 : _GEN_3068; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3070 = 8'hfe == inBytes_11 ? 8'hbb : _GEN_3069; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] outBytes_11 = 8'hff == inBytes_11 ? 8'h16 : _GEN_3070; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3073 = 8'h1 == inBytes_12 ? 8'h7c : 8'h63; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3074 = 8'h2 == inBytes_12 ? 8'h77 : _GEN_3073; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3075 = 8'h3 == inBytes_12 ? 8'h7b : _GEN_3074; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3076 = 8'h4 == inBytes_12 ? 8'hf2 : _GEN_3075; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3077 = 8'h5 == inBytes_12 ? 8'h6b : _GEN_3076; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3078 = 8'h6 == inBytes_12 ? 8'h6f : _GEN_3077; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3079 = 8'h7 == inBytes_12 ? 8'hc5 : _GEN_3078; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3080 = 8'h8 == inBytes_12 ? 8'h30 : _GEN_3079; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3081 = 8'h9 == inBytes_12 ? 8'h1 : _GEN_3080; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3082 = 8'ha == inBytes_12 ? 8'h67 : _GEN_3081; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3083 = 8'hb == inBytes_12 ? 8'h2b : _GEN_3082; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3084 = 8'hc == inBytes_12 ? 8'hfe : _GEN_3083; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3085 = 8'hd == inBytes_12 ? 8'hd7 : _GEN_3084; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3086 = 8'he == inBytes_12 ? 8'hab : _GEN_3085; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3087 = 8'hf == inBytes_12 ? 8'h76 : _GEN_3086; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3088 = 8'h10 == inBytes_12 ? 8'hca : _GEN_3087; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3089 = 8'h11 == inBytes_12 ? 8'h82 : _GEN_3088; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3090 = 8'h12 == inBytes_12 ? 8'hc9 : _GEN_3089; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3091 = 8'h13 == inBytes_12 ? 8'h7d : _GEN_3090; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3092 = 8'h14 == inBytes_12 ? 8'hfa : _GEN_3091; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3093 = 8'h15 == inBytes_12 ? 8'h59 : _GEN_3092; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3094 = 8'h16 == inBytes_12 ? 8'h47 : _GEN_3093; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3095 = 8'h17 == inBytes_12 ? 8'hf0 : _GEN_3094; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3096 = 8'h18 == inBytes_12 ? 8'had : _GEN_3095; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3097 = 8'h19 == inBytes_12 ? 8'hd4 : _GEN_3096; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3098 = 8'h1a == inBytes_12 ? 8'ha2 : _GEN_3097; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3099 = 8'h1b == inBytes_12 ? 8'haf : _GEN_3098; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3100 = 8'h1c == inBytes_12 ? 8'h9c : _GEN_3099; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3101 = 8'h1d == inBytes_12 ? 8'ha4 : _GEN_3100; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3102 = 8'h1e == inBytes_12 ? 8'h72 : _GEN_3101; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3103 = 8'h1f == inBytes_12 ? 8'hc0 : _GEN_3102; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3104 = 8'h20 == inBytes_12 ? 8'hb7 : _GEN_3103; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3105 = 8'h21 == inBytes_12 ? 8'hfd : _GEN_3104; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3106 = 8'h22 == inBytes_12 ? 8'h93 : _GEN_3105; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3107 = 8'h23 == inBytes_12 ? 8'h26 : _GEN_3106; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3108 = 8'h24 == inBytes_12 ? 8'h36 : _GEN_3107; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3109 = 8'h25 == inBytes_12 ? 8'h3f : _GEN_3108; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3110 = 8'h26 == inBytes_12 ? 8'hf7 : _GEN_3109; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3111 = 8'h27 == inBytes_12 ? 8'hcc : _GEN_3110; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3112 = 8'h28 == inBytes_12 ? 8'h34 : _GEN_3111; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3113 = 8'h29 == inBytes_12 ? 8'ha5 : _GEN_3112; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3114 = 8'h2a == inBytes_12 ? 8'he5 : _GEN_3113; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3115 = 8'h2b == inBytes_12 ? 8'hf1 : _GEN_3114; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3116 = 8'h2c == inBytes_12 ? 8'h71 : _GEN_3115; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3117 = 8'h2d == inBytes_12 ? 8'hd8 : _GEN_3116; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3118 = 8'h2e == inBytes_12 ? 8'h31 : _GEN_3117; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3119 = 8'h2f == inBytes_12 ? 8'h15 : _GEN_3118; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3120 = 8'h30 == inBytes_12 ? 8'h4 : _GEN_3119; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3121 = 8'h31 == inBytes_12 ? 8'hc7 : _GEN_3120; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3122 = 8'h32 == inBytes_12 ? 8'h23 : _GEN_3121; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3123 = 8'h33 == inBytes_12 ? 8'hc3 : _GEN_3122; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3124 = 8'h34 == inBytes_12 ? 8'h18 : _GEN_3123; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3125 = 8'h35 == inBytes_12 ? 8'h96 : _GEN_3124; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3126 = 8'h36 == inBytes_12 ? 8'h5 : _GEN_3125; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3127 = 8'h37 == inBytes_12 ? 8'h9a : _GEN_3126; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3128 = 8'h38 == inBytes_12 ? 8'h7 : _GEN_3127; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3129 = 8'h39 == inBytes_12 ? 8'h12 : _GEN_3128; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3130 = 8'h3a == inBytes_12 ? 8'h80 : _GEN_3129; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3131 = 8'h3b == inBytes_12 ? 8'he2 : _GEN_3130; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3132 = 8'h3c == inBytes_12 ? 8'heb : _GEN_3131; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3133 = 8'h3d == inBytes_12 ? 8'h27 : _GEN_3132; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3134 = 8'h3e == inBytes_12 ? 8'hb2 : _GEN_3133; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3135 = 8'h3f == inBytes_12 ? 8'h75 : _GEN_3134; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3136 = 8'h40 == inBytes_12 ? 8'h9 : _GEN_3135; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3137 = 8'h41 == inBytes_12 ? 8'h83 : _GEN_3136; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3138 = 8'h42 == inBytes_12 ? 8'h2c : _GEN_3137; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3139 = 8'h43 == inBytes_12 ? 8'h1a : _GEN_3138; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3140 = 8'h44 == inBytes_12 ? 8'h1b : _GEN_3139; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3141 = 8'h45 == inBytes_12 ? 8'h6e : _GEN_3140; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3142 = 8'h46 == inBytes_12 ? 8'h5a : _GEN_3141; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3143 = 8'h47 == inBytes_12 ? 8'ha0 : _GEN_3142; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3144 = 8'h48 == inBytes_12 ? 8'h52 : _GEN_3143; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3145 = 8'h49 == inBytes_12 ? 8'h3b : _GEN_3144; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3146 = 8'h4a == inBytes_12 ? 8'hd6 : _GEN_3145; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3147 = 8'h4b == inBytes_12 ? 8'hb3 : _GEN_3146; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3148 = 8'h4c == inBytes_12 ? 8'h29 : _GEN_3147; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3149 = 8'h4d == inBytes_12 ? 8'he3 : _GEN_3148; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3150 = 8'h4e == inBytes_12 ? 8'h2f : _GEN_3149; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3151 = 8'h4f == inBytes_12 ? 8'h84 : _GEN_3150; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3152 = 8'h50 == inBytes_12 ? 8'h53 : _GEN_3151; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3153 = 8'h51 == inBytes_12 ? 8'hd1 : _GEN_3152; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3154 = 8'h52 == inBytes_12 ? 8'h0 : _GEN_3153; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3155 = 8'h53 == inBytes_12 ? 8'hed : _GEN_3154; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3156 = 8'h54 == inBytes_12 ? 8'h20 : _GEN_3155; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3157 = 8'h55 == inBytes_12 ? 8'hfc : _GEN_3156; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3158 = 8'h56 == inBytes_12 ? 8'hb1 : _GEN_3157; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3159 = 8'h57 == inBytes_12 ? 8'h5b : _GEN_3158; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3160 = 8'h58 == inBytes_12 ? 8'h6a : _GEN_3159; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3161 = 8'h59 == inBytes_12 ? 8'hcb : _GEN_3160; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3162 = 8'h5a == inBytes_12 ? 8'hbe : _GEN_3161; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3163 = 8'h5b == inBytes_12 ? 8'h39 : _GEN_3162; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3164 = 8'h5c == inBytes_12 ? 8'h4a : _GEN_3163; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3165 = 8'h5d == inBytes_12 ? 8'h4c : _GEN_3164; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3166 = 8'h5e == inBytes_12 ? 8'h58 : _GEN_3165; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3167 = 8'h5f == inBytes_12 ? 8'hcf : _GEN_3166; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3168 = 8'h60 == inBytes_12 ? 8'hd0 : _GEN_3167; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3169 = 8'h61 == inBytes_12 ? 8'hef : _GEN_3168; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3170 = 8'h62 == inBytes_12 ? 8'haa : _GEN_3169; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3171 = 8'h63 == inBytes_12 ? 8'hfb : _GEN_3170; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3172 = 8'h64 == inBytes_12 ? 8'h43 : _GEN_3171; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3173 = 8'h65 == inBytes_12 ? 8'h4d : _GEN_3172; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3174 = 8'h66 == inBytes_12 ? 8'h33 : _GEN_3173; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3175 = 8'h67 == inBytes_12 ? 8'h85 : _GEN_3174; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3176 = 8'h68 == inBytes_12 ? 8'h45 : _GEN_3175; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3177 = 8'h69 == inBytes_12 ? 8'hf9 : _GEN_3176; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3178 = 8'h6a == inBytes_12 ? 8'h2 : _GEN_3177; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3179 = 8'h6b == inBytes_12 ? 8'h7f : _GEN_3178; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3180 = 8'h6c == inBytes_12 ? 8'h50 : _GEN_3179; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3181 = 8'h6d == inBytes_12 ? 8'h3c : _GEN_3180; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3182 = 8'h6e == inBytes_12 ? 8'h9f : _GEN_3181; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3183 = 8'h6f == inBytes_12 ? 8'ha8 : _GEN_3182; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3184 = 8'h70 == inBytes_12 ? 8'h51 : _GEN_3183; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3185 = 8'h71 == inBytes_12 ? 8'ha3 : _GEN_3184; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3186 = 8'h72 == inBytes_12 ? 8'h40 : _GEN_3185; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3187 = 8'h73 == inBytes_12 ? 8'h8f : _GEN_3186; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3188 = 8'h74 == inBytes_12 ? 8'h92 : _GEN_3187; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3189 = 8'h75 == inBytes_12 ? 8'h9d : _GEN_3188; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3190 = 8'h76 == inBytes_12 ? 8'h38 : _GEN_3189; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3191 = 8'h77 == inBytes_12 ? 8'hf5 : _GEN_3190; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3192 = 8'h78 == inBytes_12 ? 8'hbc : _GEN_3191; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3193 = 8'h79 == inBytes_12 ? 8'hb6 : _GEN_3192; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3194 = 8'h7a == inBytes_12 ? 8'hda : _GEN_3193; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3195 = 8'h7b == inBytes_12 ? 8'h21 : _GEN_3194; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3196 = 8'h7c == inBytes_12 ? 8'h10 : _GEN_3195; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3197 = 8'h7d == inBytes_12 ? 8'hff : _GEN_3196; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3198 = 8'h7e == inBytes_12 ? 8'hf3 : _GEN_3197; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3199 = 8'h7f == inBytes_12 ? 8'hd2 : _GEN_3198; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3200 = 8'h80 == inBytes_12 ? 8'hcd : _GEN_3199; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3201 = 8'h81 == inBytes_12 ? 8'hc : _GEN_3200; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3202 = 8'h82 == inBytes_12 ? 8'h13 : _GEN_3201; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3203 = 8'h83 == inBytes_12 ? 8'hec : _GEN_3202; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3204 = 8'h84 == inBytes_12 ? 8'h5f : _GEN_3203; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3205 = 8'h85 == inBytes_12 ? 8'h97 : _GEN_3204; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3206 = 8'h86 == inBytes_12 ? 8'h44 : _GEN_3205; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3207 = 8'h87 == inBytes_12 ? 8'h17 : _GEN_3206; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3208 = 8'h88 == inBytes_12 ? 8'hc4 : _GEN_3207; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3209 = 8'h89 == inBytes_12 ? 8'ha7 : _GEN_3208; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3210 = 8'h8a == inBytes_12 ? 8'h7e : _GEN_3209; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3211 = 8'h8b == inBytes_12 ? 8'h3d : _GEN_3210; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3212 = 8'h8c == inBytes_12 ? 8'h64 : _GEN_3211; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3213 = 8'h8d == inBytes_12 ? 8'h5d : _GEN_3212; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3214 = 8'h8e == inBytes_12 ? 8'h19 : _GEN_3213; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3215 = 8'h8f == inBytes_12 ? 8'h73 : _GEN_3214; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3216 = 8'h90 == inBytes_12 ? 8'h60 : _GEN_3215; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3217 = 8'h91 == inBytes_12 ? 8'h81 : _GEN_3216; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3218 = 8'h92 == inBytes_12 ? 8'h4f : _GEN_3217; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3219 = 8'h93 == inBytes_12 ? 8'hdc : _GEN_3218; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3220 = 8'h94 == inBytes_12 ? 8'h22 : _GEN_3219; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3221 = 8'h95 == inBytes_12 ? 8'h2a : _GEN_3220; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3222 = 8'h96 == inBytes_12 ? 8'h90 : _GEN_3221; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3223 = 8'h97 == inBytes_12 ? 8'h88 : _GEN_3222; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3224 = 8'h98 == inBytes_12 ? 8'h46 : _GEN_3223; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3225 = 8'h99 == inBytes_12 ? 8'hee : _GEN_3224; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3226 = 8'h9a == inBytes_12 ? 8'hb8 : _GEN_3225; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3227 = 8'h9b == inBytes_12 ? 8'h14 : _GEN_3226; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3228 = 8'h9c == inBytes_12 ? 8'hde : _GEN_3227; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3229 = 8'h9d == inBytes_12 ? 8'h5e : _GEN_3228; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3230 = 8'h9e == inBytes_12 ? 8'hb : _GEN_3229; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3231 = 8'h9f == inBytes_12 ? 8'hdb : _GEN_3230; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3232 = 8'ha0 == inBytes_12 ? 8'he0 : _GEN_3231; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3233 = 8'ha1 == inBytes_12 ? 8'h32 : _GEN_3232; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3234 = 8'ha2 == inBytes_12 ? 8'h3a : _GEN_3233; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3235 = 8'ha3 == inBytes_12 ? 8'ha : _GEN_3234; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3236 = 8'ha4 == inBytes_12 ? 8'h49 : _GEN_3235; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3237 = 8'ha5 == inBytes_12 ? 8'h6 : _GEN_3236; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3238 = 8'ha6 == inBytes_12 ? 8'h24 : _GEN_3237; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3239 = 8'ha7 == inBytes_12 ? 8'h5c : _GEN_3238; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3240 = 8'ha8 == inBytes_12 ? 8'hc2 : _GEN_3239; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3241 = 8'ha9 == inBytes_12 ? 8'hd3 : _GEN_3240; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3242 = 8'haa == inBytes_12 ? 8'hac : _GEN_3241; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3243 = 8'hab == inBytes_12 ? 8'h62 : _GEN_3242; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3244 = 8'hac == inBytes_12 ? 8'h91 : _GEN_3243; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3245 = 8'had == inBytes_12 ? 8'h95 : _GEN_3244; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3246 = 8'hae == inBytes_12 ? 8'he4 : _GEN_3245; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3247 = 8'haf == inBytes_12 ? 8'h79 : _GEN_3246; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3248 = 8'hb0 == inBytes_12 ? 8'he7 : _GEN_3247; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3249 = 8'hb1 == inBytes_12 ? 8'hc8 : _GEN_3248; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3250 = 8'hb2 == inBytes_12 ? 8'h37 : _GEN_3249; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3251 = 8'hb3 == inBytes_12 ? 8'h6d : _GEN_3250; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3252 = 8'hb4 == inBytes_12 ? 8'h8d : _GEN_3251; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3253 = 8'hb5 == inBytes_12 ? 8'hd5 : _GEN_3252; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3254 = 8'hb6 == inBytes_12 ? 8'h4e : _GEN_3253; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3255 = 8'hb7 == inBytes_12 ? 8'ha9 : _GEN_3254; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3256 = 8'hb8 == inBytes_12 ? 8'h6c : _GEN_3255; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3257 = 8'hb9 == inBytes_12 ? 8'h56 : _GEN_3256; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3258 = 8'hba == inBytes_12 ? 8'hf4 : _GEN_3257; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3259 = 8'hbb == inBytes_12 ? 8'hea : _GEN_3258; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3260 = 8'hbc == inBytes_12 ? 8'h65 : _GEN_3259; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3261 = 8'hbd == inBytes_12 ? 8'h7a : _GEN_3260; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3262 = 8'hbe == inBytes_12 ? 8'hae : _GEN_3261; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3263 = 8'hbf == inBytes_12 ? 8'h8 : _GEN_3262; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3264 = 8'hc0 == inBytes_12 ? 8'hba : _GEN_3263; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3265 = 8'hc1 == inBytes_12 ? 8'h78 : _GEN_3264; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3266 = 8'hc2 == inBytes_12 ? 8'h25 : _GEN_3265; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3267 = 8'hc3 == inBytes_12 ? 8'h2e : _GEN_3266; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3268 = 8'hc4 == inBytes_12 ? 8'h1c : _GEN_3267; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3269 = 8'hc5 == inBytes_12 ? 8'ha6 : _GEN_3268; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3270 = 8'hc6 == inBytes_12 ? 8'hb4 : _GEN_3269; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3271 = 8'hc7 == inBytes_12 ? 8'hc6 : _GEN_3270; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3272 = 8'hc8 == inBytes_12 ? 8'he8 : _GEN_3271; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3273 = 8'hc9 == inBytes_12 ? 8'hdd : _GEN_3272; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3274 = 8'hca == inBytes_12 ? 8'h74 : _GEN_3273; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3275 = 8'hcb == inBytes_12 ? 8'h1f : _GEN_3274; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3276 = 8'hcc == inBytes_12 ? 8'h4b : _GEN_3275; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3277 = 8'hcd == inBytes_12 ? 8'hbd : _GEN_3276; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3278 = 8'hce == inBytes_12 ? 8'h8b : _GEN_3277; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3279 = 8'hcf == inBytes_12 ? 8'h8a : _GEN_3278; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3280 = 8'hd0 == inBytes_12 ? 8'h70 : _GEN_3279; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3281 = 8'hd1 == inBytes_12 ? 8'h3e : _GEN_3280; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3282 = 8'hd2 == inBytes_12 ? 8'hb5 : _GEN_3281; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3283 = 8'hd3 == inBytes_12 ? 8'h66 : _GEN_3282; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3284 = 8'hd4 == inBytes_12 ? 8'h48 : _GEN_3283; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3285 = 8'hd5 == inBytes_12 ? 8'h3 : _GEN_3284; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3286 = 8'hd6 == inBytes_12 ? 8'hf6 : _GEN_3285; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3287 = 8'hd7 == inBytes_12 ? 8'he : _GEN_3286; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3288 = 8'hd8 == inBytes_12 ? 8'h61 : _GEN_3287; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3289 = 8'hd9 == inBytes_12 ? 8'h35 : _GEN_3288; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3290 = 8'hda == inBytes_12 ? 8'h57 : _GEN_3289; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3291 = 8'hdb == inBytes_12 ? 8'hb9 : _GEN_3290; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3292 = 8'hdc == inBytes_12 ? 8'h86 : _GEN_3291; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3293 = 8'hdd == inBytes_12 ? 8'hc1 : _GEN_3292; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3294 = 8'hde == inBytes_12 ? 8'h1d : _GEN_3293; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3295 = 8'hdf == inBytes_12 ? 8'h9e : _GEN_3294; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3296 = 8'he0 == inBytes_12 ? 8'he1 : _GEN_3295; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3297 = 8'he1 == inBytes_12 ? 8'hf8 : _GEN_3296; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3298 = 8'he2 == inBytes_12 ? 8'h98 : _GEN_3297; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3299 = 8'he3 == inBytes_12 ? 8'h11 : _GEN_3298; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3300 = 8'he4 == inBytes_12 ? 8'h69 : _GEN_3299; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3301 = 8'he5 == inBytes_12 ? 8'hd9 : _GEN_3300; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3302 = 8'he6 == inBytes_12 ? 8'h8e : _GEN_3301; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3303 = 8'he7 == inBytes_12 ? 8'h94 : _GEN_3302; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3304 = 8'he8 == inBytes_12 ? 8'h9b : _GEN_3303; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3305 = 8'he9 == inBytes_12 ? 8'h1e : _GEN_3304; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3306 = 8'hea == inBytes_12 ? 8'h87 : _GEN_3305; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3307 = 8'heb == inBytes_12 ? 8'he9 : _GEN_3306; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3308 = 8'hec == inBytes_12 ? 8'hce : _GEN_3307; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3309 = 8'hed == inBytes_12 ? 8'h55 : _GEN_3308; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3310 = 8'hee == inBytes_12 ? 8'h28 : _GEN_3309; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3311 = 8'hef == inBytes_12 ? 8'hdf : _GEN_3310; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3312 = 8'hf0 == inBytes_12 ? 8'h8c : _GEN_3311; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3313 = 8'hf1 == inBytes_12 ? 8'ha1 : _GEN_3312; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3314 = 8'hf2 == inBytes_12 ? 8'h89 : _GEN_3313; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3315 = 8'hf3 == inBytes_12 ? 8'hd : _GEN_3314; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3316 = 8'hf4 == inBytes_12 ? 8'hbf : _GEN_3315; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3317 = 8'hf5 == inBytes_12 ? 8'he6 : _GEN_3316; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3318 = 8'hf6 == inBytes_12 ? 8'h42 : _GEN_3317; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3319 = 8'hf7 == inBytes_12 ? 8'h68 : _GEN_3318; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3320 = 8'hf8 == inBytes_12 ? 8'h41 : _GEN_3319; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3321 = 8'hf9 == inBytes_12 ? 8'h99 : _GEN_3320; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3322 = 8'hfa == inBytes_12 ? 8'h2d : _GEN_3321; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3323 = 8'hfb == inBytes_12 ? 8'hf : _GEN_3322; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3324 = 8'hfc == inBytes_12 ? 8'hb0 : _GEN_3323; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3325 = 8'hfd == inBytes_12 ? 8'h54 : _GEN_3324; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3326 = 8'hfe == inBytes_12 ? 8'hbb : _GEN_3325; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] outBytes_12 = 8'hff == inBytes_12 ? 8'h16 : _GEN_3326; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3329 = 8'h1 == inBytes_13 ? 8'h7c : 8'h63; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3330 = 8'h2 == inBytes_13 ? 8'h77 : _GEN_3329; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3331 = 8'h3 == inBytes_13 ? 8'h7b : _GEN_3330; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3332 = 8'h4 == inBytes_13 ? 8'hf2 : _GEN_3331; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3333 = 8'h5 == inBytes_13 ? 8'h6b : _GEN_3332; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3334 = 8'h6 == inBytes_13 ? 8'h6f : _GEN_3333; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3335 = 8'h7 == inBytes_13 ? 8'hc5 : _GEN_3334; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3336 = 8'h8 == inBytes_13 ? 8'h30 : _GEN_3335; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3337 = 8'h9 == inBytes_13 ? 8'h1 : _GEN_3336; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3338 = 8'ha == inBytes_13 ? 8'h67 : _GEN_3337; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3339 = 8'hb == inBytes_13 ? 8'h2b : _GEN_3338; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3340 = 8'hc == inBytes_13 ? 8'hfe : _GEN_3339; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3341 = 8'hd == inBytes_13 ? 8'hd7 : _GEN_3340; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3342 = 8'he == inBytes_13 ? 8'hab : _GEN_3341; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3343 = 8'hf == inBytes_13 ? 8'h76 : _GEN_3342; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3344 = 8'h10 == inBytes_13 ? 8'hca : _GEN_3343; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3345 = 8'h11 == inBytes_13 ? 8'h82 : _GEN_3344; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3346 = 8'h12 == inBytes_13 ? 8'hc9 : _GEN_3345; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3347 = 8'h13 == inBytes_13 ? 8'h7d : _GEN_3346; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3348 = 8'h14 == inBytes_13 ? 8'hfa : _GEN_3347; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3349 = 8'h15 == inBytes_13 ? 8'h59 : _GEN_3348; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3350 = 8'h16 == inBytes_13 ? 8'h47 : _GEN_3349; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3351 = 8'h17 == inBytes_13 ? 8'hf0 : _GEN_3350; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3352 = 8'h18 == inBytes_13 ? 8'had : _GEN_3351; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3353 = 8'h19 == inBytes_13 ? 8'hd4 : _GEN_3352; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3354 = 8'h1a == inBytes_13 ? 8'ha2 : _GEN_3353; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3355 = 8'h1b == inBytes_13 ? 8'haf : _GEN_3354; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3356 = 8'h1c == inBytes_13 ? 8'h9c : _GEN_3355; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3357 = 8'h1d == inBytes_13 ? 8'ha4 : _GEN_3356; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3358 = 8'h1e == inBytes_13 ? 8'h72 : _GEN_3357; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3359 = 8'h1f == inBytes_13 ? 8'hc0 : _GEN_3358; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3360 = 8'h20 == inBytes_13 ? 8'hb7 : _GEN_3359; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3361 = 8'h21 == inBytes_13 ? 8'hfd : _GEN_3360; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3362 = 8'h22 == inBytes_13 ? 8'h93 : _GEN_3361; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3363 = 8'h23 == inBytes_13 ? 8'h26 : _GEN_3362; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3364 = 8'h24 == inBytes_13 ? 8'h36 : _GEN_3363; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3365 = 8'h25 == inBytes_13 ? 8'h3f : _GEN_3364; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3366 = 8'h26 == inBytes_13 ? 8'hf7 : _GEN_3365; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3367 = 8'h27 == inBytes_13 ? 8'hcc : _GEN_3366; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3368 = 8'h28 == inBytes_13 ? 8'h34 : _GEN_3367; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3369 = 8'h29 == inBytes_13 ? 8'ha5 : _GEN_3368; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3370 = 8'h2a == inBytes_13 ? 8'he5 : _GEN_3369; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3371 = 8'h2b == inBytes_13 ? 8'hf1 : _GEN_3370; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3372 = 8'h2c == inBytes_13 ? 8'h71 : _GEN_3371; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3373 = 8'h2d == inBytes_13 ? 8'hd8 : _GEN_3372; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3374 = 8'h2e == inBytes_13 ? 8'h31 : _GEN_3373; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3375 = 8'h2f == inBytes_13 ? 8'h15 : _GEN_3374; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3376 = 8'h30 == inBytes_13 ? 8'h4 : _GEN_3375; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3377 = 8'h31 == inBytes_13 ? 8'hc7 : _GEN_3376; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3378 = 8'h32 == inBytes_13 ? 8'h23 : _GEN_3377; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3379 = 8'h33 == inBytes_13 ? 8'hc3 : _GEN_3378; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3380 = 8'h34 == inBytes_13 ? 8'h18 : _GEN_3379; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3381 = 8'h35 == inBytes_13 ? 8'h96 : _GEN_3380; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3382 = 8'h36 == inBytes_13 ? 8'h5 : _GEN_3381; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3383 = 8'h37 == inBytes_13 ? 8'h9a : _GEN_3382; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3384 = 8'h38 == inBytes_13 ? 8'h7 : _GEN_3383; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3385 = 8'h39 == inBytes_13 ? 8'h12 : _GEN_3384; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3386 = 8'h3a == inBytes_13 ? 8'h80 : _GEN_3385; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3387 = 8'h3b == inBytes_13 ? 8'he2 : _GEN_3386; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3388 = 8'h3c == inBytes_13 ? 8'heb : _GEN_3387; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3389 = 8'h3d == inBytes_13 ? 8'h27 : _GEN_3388; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3390 = 8'h3e == inBytes_13 ? 8'hb2 : _GEN_3389; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3391 = 8'h3f == inBytes_13 ? 8'h75 : _GEN_3390; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3392 = 8'h40 == inBytes_13 ? 8'h9 : _GEN_3391; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3393 = 8'h41 == inBytes_13 ? 8'h83 : _GEN_3392; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3394 = 8'h42 == inBytes_13 ? 8'h2c : _GEN_3393; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3395 = 8'h43 == inBytes_13 ? 8'h1a : _GEN_3394; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3396 = 8'h44 == inBytes_13 ? 8'h1b : _GEN_3395; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3397 = 8'h45 == inBytes_13 ? 8'h6e : _GEN_3396; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3398 = 8'h46 == inBytes_13 ? 8'h5a : _GEN_3397; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3399 = 8'h47 == inBytes_13 ? 8'ha0 : _GEN_3398; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3400 = 8'h48 == inBytes_13 ? 8'h52 : _GEN_3399; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3401 = 8'h49 == inBytes_13 ? 8'h3b : _GEN_3400; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3402 = 8'h4a == inBytes_13 ? 8'hd6 : _GEN_3401; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3403 = 8'h4b == inBytes_13 ? 8'hb3 : _GEN_3402; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3404 = 8'h4c == inBytes_13 ? 8'h29 : _GEN_3403; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3405 = 8'h4d == inBytes_13 ? 8'he3 : _GEN_3404; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3406 = 8'h4e == inBytes_13 ? 8'h2f : _GEN_3405; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3407 = 8'h4f == inBytes_13 ? 8'h84 : _GEN_3406; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3408 = 8'h50 == inBytes_13 ? 8'h53 : _GEN_3407; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3409 = 8'h51 == inBytes_13 ? 8'hd1 : _GEN_3408; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3410 = 8'h52 == inBytes_13 ? 8'h0 : _GEN_3409; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3411 = 8'h53 == inBytes_13 ? 8'hed : _GEN_3410; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3412 = 8'h54 == inBytes_13 ? 8'h20 : _GEN_3411; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3413 = 8'h55 == inBytes_13 ? 8'hfc : _GEN_3412; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3414 = 8'h56 == inBytes_13 ? 8'hb1 : _GEN_3413; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3415 = 8'h57 == inBytes_13 ? 8'h5b : _GEN_3414; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3416 = 8'h58 == inBytes_13 ? 8'h6a : _GEN_3415; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3417 = 8'h59 == inBytes_13 ? 8'hcb : _GEN_3416; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3418 = 8'h5a == inBytes_13 ? 8'hbe : _GEN_3417; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3419 = 8'h5b == inBytes_13 ? 8'h39 : _GEN_3418; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3420 = 8'h5c == inBytes_13 ? 8'h4a : _GEN_3419; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3421 = 8'h5d == inBytes_13 ? 8'h4c : _GEN_3420; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3422 = 8'h5e == inBytes_13 ? 8'h58 : _GEN_3421; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3423 = 8'h5f == inBytes_13 ? 8'hcf : _GEN_3422; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3424 = 8'h60 == inBytes_13 ? 8'hd0 : _GEN_3423; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3425 = 8'h61 == inBytes_13 ? 8'hef : _GEN_3424; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3426 = 8'h62 == inBytes_13 ? 8'haa : _GEN_3425; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3427 = 8'h63 == inBytes_13 ? 8'hfb : _GEN_3426; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3428 = 8'h64 == inBytes_13 ? 8'h43 : _GEN_3427; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3429 = 8'h65 == inBytes_13 ? 8'h4d : _GEN_3428; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3430 = 8'h66 == inBytes_13 ? 8'h33 : _GEN_3429; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3431 = 8'h67 == inBytes_13 ? 8'h85 : _GEN_3430; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3432 = 8'h68 == inBytes_13 ? 8'h45 : _GEN_3431; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3433 = 8'h69 == inBytes_13 ? 8'hf9 : _GEN_3432; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3434 = 8'h6a == inBytes_13 ? 8'h2 : _GEN_3433; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3435 = 8'h6b == inBytes_13 ? 8'h7f : _GEN_3434; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3436 = 8'h6c == inBytes_13 ? 8'h50 : _GEN_3435; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3437 = 8'h6d == inBytes_13 ? 8'h3c : _GEN_3436; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3438 = 8'h6e == inBytes_13 ? 8'h9f : _GEN_3437; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3439 = 8'h6f == inBytes_13 ? 8'ha8 : _GEN_3438; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3440 = 8'h70 == inBytes_13 ? 8'h51 : _GEN_3439; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3441 = 8'h71 == inBytes_13 ? 8'ha3 : _GEN_3440; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3442 = 8'h72 == inBytes_13 ? 8'h40 : _GEN_3441; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3443 = 8'h73 == inBytes_13 ? 8'h8f : _GEN_3442; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3444 = 8'h74 == inBytes_13 ? 8'h92 : _GEN_3443; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3445 = 8'h75 == inBytes_13 ? 8'h9d : _GEN_3444; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3446 = 8'h76 == inBytes_13 ? 8'h38 : _GEN_3445; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3447 = 8'h77 == inBytes_13 ? 8'hf5 : _GEN_3446; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3448 = 8'h78 == inBytes_13 ? 8'hbc : _GEN_3447; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3449 = 8'h79 == inBytes_13 ? 8'hb6 : _GEN_3448; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3450 = 8'h7a == inBytes_13 ? 8'hda : _GEN_3449; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3451 = 8'h7b == inBytes_13 ? 8'h21 : _GEN_3450; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3452 = 8'h7c == inBytes_13 ? 8'h10 : _GEN_3451; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3453 = 8'h7d == inBytes_13 ? 8'hff : _GEN_3452; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3454 = 8'h7e == inBytes_13 ? 8'hf3 : _GEN_3453; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3455 = 8'h7f == inBytes_13 ? 8'hd2 : _GEN_3454; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3456 = 8'h80 == inBytes_13 ? 8'hcd : _GEN_3455; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3457 = 8'h81 == inBytes_13 ? 8'hc : _GEN_3456; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3458 = 8'h82 == inBytes_13 ? 8'h13 : _GEN_3457; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3459 = 8'h83 == inBytes_13 ? 8'hec : _GEN_3458; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3460 = 8'h84 == inBytes_13 ? 8'h5f : _GEN_3459; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3461 = 8'h85 == inBytes_13 ? 8'h97 : _GEN_3460; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3462 = 8'h86 == inBytes_13 ? 8'h44 : _GEN_3461; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3463 = 8'h87 == inBytes_13 ? 8'h17 : _GEN_3462; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3464 = 8'h88 == inBytes_13 ? 8'hc4 : _GEN_3463; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3465 = 8'h89 == inBytes_13 ? 8'ha7 : _GEN_3464; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3466 = 8'h8a == inBytes_13 ? 8'h7e : _GEN_3465; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3467 = 8'h8b == inBytes_13 ? 8'h3d : _GEN_3466; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3468 = 8'h8c == inBytes_13 ? 8'h64 : _GEN_3467; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3469 = 8'h8d == inBytes_13 ? 8'h5d : _GEN_3468; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3470 = 8'h8e == inBytes_13 ? 8'h19 : _GEN_3469; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3471 = 8'h8f == inBytes_13 ? 8'h73 : _GEN_3470; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3472 = 8'h90 == inBytes_13 ? 8'h60 : _GEN_3471; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3473 = 8'h91 == inBytes_13 ? 8'h81 : _GEN_3472; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3474 = 8'h92 == inBytes_13 ? 8'h4f : _GEN_3473; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3475 = 8'h93 == inBytes_13 ? 8'hdc : _GEN_3474; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3476 = 8'h94 == inBytes_13 ? 8'h22 : _GEN_3475; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3477 = 8'h95 == inBytes_13 ? 8'h2a : _GEN_3476; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3478 = 8'h96 == inBytes_13 ? 8'h90 : _GEN_3477; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3479 = 8'h97 == inBytes_13 ? 8'h88 : _GEN_3478; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3480 = 8'h98 == inBytes_13 ? 8'h46 : _GEN_3479; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3481 = 8'h99 == inBytes_13 ? 8'hee : _GEN_3480; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3482 = 8'h9a == inBytes_13 ? 8'hb8 : _GEN_3481; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3483 = 8'h9b == inBytes_13 ? 8'h14 : _GEN_3482; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3484 = 8'h9c == inBytes_13 ? 8'hde : _GEN_3483; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3485 = 8'h9d == inBytes_13 ? 8'h5e : _GEN_3484; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3486 = 8'h9e == inBytes_13 ? 8'hb : _GEN_3485; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3487 = 8'h9f == inBytes_13 ? 8'hdb : _GEN_3486; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3488 = 8'ha0 == inBytes_13 ? 8'he0 : _GEN_3487; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3489 = 8'ha1 == inBytes_13 ? 8'h32 : _GEN_3488; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3490 = 8'ha2 == inBytes_13 ? 8'h3a : _GEN_3489; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3491 = 8'ha3 == inBytes_13 ? 8'ha : _GEN_3490; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3492 = 8'ha4 == inBytes_13 ? 8'h49 : _GEN_3491; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3493 = 8'ha5 == inBytes_13 ? 8'h6 : _GEN_3492; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3494 = 8'ha6 == inBytes_13 ? 8'h24 : _GEN_3493; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3495 = 8'ha7 == inBytes_13 ? 8'h5c : _GEN_3494; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3496 = 8'ha8 == inBytes_13 ? 8'hc2 : _GEN_3495; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3497 = 8'ha9 == inBytes_13 ? 8'hd3 : _GEN_3496; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3498 = 8'haa == inBytes_13 ? 8'hac : _GEN_3497; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3499 = 8'hab == inBytes_13 ? 8'h62 : _GEN_3498; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3500 = 8'hac == inBytes_13 ? 8'h91 : _GEN_3499; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3501 = 8'had == inBytes_13 ? 8'h95 : _GEN_3500; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3502 = 8'hae == inBytes_13 ? 8'he4 : _GEN_3501; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3503 = 8'haf == inBytes_13 ? 8'h79 : _GEN_3502; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3504 = 8'hb0 == inBytes_13 ? 8'he7 : _GEN_3503; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3505 = 8'hb1 == inBytes_13 ? 8'hc8 : _GEN_3504; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3506 = 8'hb2 == inBytes_13 ? 8'h37 : _GEN_3505; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3507 = 8'hb3 == inBytes_13 ? 8'h6d : _GEN_3506; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3508 = 8'hb4 == inBytes_13 ? 8'h8d : _GEN_3507; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3509 = 8'hb5 == inBytes_13 ? 8'hd5 : _GEN_3508; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3510 = 8'hb6 == inBytes_13 ? 8'h4e : _GEN_3509; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3511 = 8'hb7 == inBytes_13 ? 8'ha9 : _GEN_3510; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3512 = 8'hb8 == inBytes_13 ? 8'h6c : _GEN_3511; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3513 = 8'hb9 == inBytes_13 ? 8'h56 : _GEN_3512; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3514 = 8'hba == inBytes_13 ? 8'hf4 : _GEN_3513; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3515 = 8'hbb == inBytes_13 ? 8'hea : _GEN_3514; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3516 = 8'hbc == inBytes_13 ? 8'h65 : _GEN_3515; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3517 = 8'hbd == inBytes_13 ? 8'h7a : _GEN_3516; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3518 = 8'hbe == inBytes_13 ? 8'hae : _GEN_3517; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3519 = 8'hbf == inBytes_13 ? 8'h8 : _GEN_3518; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3520 = 8'hc0 == inBytes_13 ? 8'hba : _GEN_3519; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3521 = 8'hc1 == inBytes_13 ? 8'h78 : _GEN_3520; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3522 = 8'hc2 == inBytes_13 ? 8'h25 : _GEN_3521; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3523 = 8'hc3 == inBytes_13 ? 8'h2e : _GEN_3522; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3524 = 8'hc4 == inBytes_13 ? 8'h1c : _GEN_3523; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3525 = 8'hc5 == inBytes_13 ? 8'ha6 : _GEN_3524; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3526 = 8'hc6 == inBytes_13 ? 8'hb4 : _GEN_3525; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3527 = 8'hc7 == inBytes_13 ? 8'hc6 : _GEN_3526; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3528 = 8'hc8 == inBytes_13 ? 8'he8 : _GEN_3527; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3529 = 8'hc9 == inBytes_13 ? 8'hdd : _GEN_3528; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3530 = 8'hca == inBytes_13 ? 8'h74 : _GEN_3529; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3531 = 8'hcb == inBytes_13 ? 8'h1f : _GEN_3530; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3532 = 8'hcc == inBytes_13 ? 8'h4b : _GEN_3531; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3533 = 8'hcd == inBytes_13 ? 8'hbd : _GEN_3532; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3534 = 8'hce == inBytes_13 ? 8'h8b : _GEN_3533; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3535 = 8'hcf == inBytes_13 ? 8'h8a : _GEN_3534; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3536 = 8'hd0 == inBytes_13 ? 8'h70 : _GEN_3535; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3537 = 8'hd1 == inBytes_13 ? 8'h3e : _GEN_3536; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3538 = 8'hd2 == inBytes_13 ? 8'hb5 : _GEN_3537; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3539 = 8'hd3 == inBytes_13 ? 8'h66 : _GEN_3538; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3540 = 8'hd4 == inBytes_13 ? 8'h48 : _GEN_3539; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3541 = 8'hd5 == inBytes_13 ? 8'h3 : _GEN_3540; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3542 = 8'hd6 == inBytes_13 ? 8'hf6 : _GEN_3541; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3543 = 8'hd7 == inBytes_13 ? 8'he : _GEN_3542; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3544 = 8'hd8 == inBytes_13 ? 8'h61 : _GEN_3543; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3545 = 8'hd9 == inBytes_13 ? 8'h35 : _GEN_3544; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3546 = 8'hda == inBytes_13 ? 8'h57 : _GEN_3545; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3547 = 8'hdb == inBytes_13 ? 8'hb9 : _GEN_3546; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3548 = 8'hdc == inBytes_13 ? 8'h86 : _GEN_3547; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3549 = 8'hdd == inBytes_13 ? 8'hc1 : _GEN_3548; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3550 = 8'hde == inBytes_13 ? 8'h1d : _GEN_3549; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3551 = 8'hdf == inBytes_13 ? 8'h9e : _GEN_3550; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3552 = 8'he0 == inBytes_13 ? 8'he1 : _GEN_3551; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3553 = 8'he1 == inBytes_13 ? 8'hf8 : _GEN_3552; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3554 = 8'he2 == inBytes_13 ? 8'h98 : _GEN_3553; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3555 = 8'he3 == inBytes_13 ? 8'h11 : _GEN_3554; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3556 = 8'he4 == inBytes_13 ? 8'h69 : _GEN_3555; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3557 = 8'he5 == inBytes_13 ? 8'hd9 : _GEN_3556; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3558 = 8'he6 == inBytes_13 ? 8'h8e : _GEN_3557; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3559 = 8'he7 == inBytes_13 ? 8'h94 : _GEN_3558; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3560 = 8'he8 == inBytes_13 ? 8'h9b : _GEN_3559; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3561 = 8'he9 == inBytes_13 ? 8'h1e : _GEN_3560; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3562 = 8'hea == inBytes_13 ? 8'h87 : _GEN_3561; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3563 = 8'heb == inBytes_13 ? 8'he9 : _GEN_3562; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3564 = 8'hec == inBytes_13 ? 8'hce : _GEN_3563; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3565 = 8'hed == inBytes_13 ? 8'h55 : _GEN_3564; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3566 = 8'hee == inBytes_13 ? 8'h28 : _GEN_3565; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3567 = 8'hef == inBytes_13 ? 8'hdf : _GEN_3566; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3568 = 8'hf0 == inBytes_13 ? 8'h8c : _GEN_3567; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3569 = 8'hf1 == inBytes_13 ? 8'ha1 : _GEN_3568; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3570 = 8'hf2 == inBytes_13 ? 8'h89 : _GEN_3569; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3571 = 8'hf3 == inBytes_13 ? 8'hd : _GEN_3570; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3572 = 8'hf4 == inBytes_13 ? 8'hbf : _GEN_3571; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3573 = 8'hf5 == inBytes_13 ? 8'he6 : _GEN_3572; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3574 = 8'hf6 == inBytes_13 ? 8'h42 : _GEN_3573; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3575 = 8'hf7 == inBytes_13 ? 8'h68 : _GEN_3574; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3576 = 8'hf8 == inBytes_13 ? 8'h41 : _GEN_3575; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3577 = 8'hf9 == inBytes_13 ? 8'h99 : _GEN_3576; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3578 = 8'hfa == inBytes_13 ? 8'h2d : _GEN_3577; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3579 = 8'hfb == inBytes_13 ? 8'hf : _GEN_3578; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3580 = 8'hfc == inBytes_13 ? 8'hb0 : _GEN_3579; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3581 = 8'hfd == inBytes_13 ? 8'h54 : _GEN_3580; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3582 = 8'hfe == inBytes_13 ? 8'hbb : _GEN_3581; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] outBytes_13 = 8'hff == inBytes_13 ? 8'h16 : _GEN_3582; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3585 = 8'h1 == inBytes_14 ? 8'h7c : 8'h63; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3586 = 8'h2 == inBytes_14 ? 8'h77 : _GEN_3585; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3587 = 8'h3 == inBytes_14 ? 8'h7b : _GEN_3586; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3588 = 8'h4 == inBytes_14 ? 8'hf2 : _GEN_3587; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3589 = 8'h5 == inBytes_14 ? 8'h6b : _GEN_3588; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3590 = 8'h6 == inBytes_14 ? 8'h6f : _GEN_3589; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3591 = 8'h7 == inBytes_14 ? 8'hc5 : _GEN_3590; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3592 = 8'h8 == inBytes_14 ? 8'h30 : _GEN_3591; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3593 = 8'h9 == inBytes_14 ? 8'h1 : _GEN_3592; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3594 = 8'ha == inBytes_14 ? 8'h67 : _GEN_3593; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3595 = 8'hb == inBytes_14 ? 8'h2b : _GEN_3594; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3596 = 8'hc == inBytes_14 ? 8'hfe : _GEN_3595; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3597 = 8'hd == inBytes_14 ? 8'hd7 : _GEN_3596; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3598 = 8'he == inBytes_14 ? 8'hab : _GEN_3597; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3599 = 8'hf == inBytes_14 ? 8'h76 : _GEN_3598; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3600 = 8'h10 == inBytes_14 ? 8'hca : _GEN_3599; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3601 = 8'h11 == inBytes_14 ? 8'h82 : _GEN_3600; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3602 = 8'h12 == inBytes_14 ? 8'hc9 : _GEN_3601; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3603 = 8'h13 == inBytes_14 ? 8'h7d : _GEN_3602; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3604 = 8'h14 == inBytes_14 ? 8'hfa : _GEN_3603; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3605 = 8'h15 == inBytes_14 ? 8'h59 : _GEN_3604; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3606 = 8'h16 == inBytes_14 ? 8'h47 : _GEN_3605; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3607 = 8'h17 == inBytes_14 ? 8'hf0 : _GEN_3606; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3608 = 8'h18 == inBytes_14 ? 8'had : _GEN_3607; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3609 = 8'h19 == inBytes_14 ? 8'hd4 : _GEN_3608; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3610 = 8'h1a == inBytes_14 ? 8'ha2 : _GEN_3609; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3611 = 8'h1b == inBytes_14 ? 8'haf : _GEN_3610; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3612 = 8'h1c == inBytes_14 ? 8'h9c : _GEN_3611; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3613 = 8'h1d == inBytes_14 ? 8'ha4 : _GEN_3612; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3614 = 8'h1e == inBytes_14 ? 8'h72 : _GEN_3613; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3615 = 8'h1f == inBytes_14 ? 8'hc0 : _GEN_3614; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3616 = 8'h20 == inBytes_14 ? 8'hb7 : _GEN_3615; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3617 = 8'h21 == inBytes_14 ? 8'hfd : _GEN_3616; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3618 = 8'h22 == inBytes_14 ? 8'h93 : _GEN_3617; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3619 = 8'h23 == inBytes_14 ? 8'h26 : _GEN_3618; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3620 = 8'h24 == inBytes_14 ? 8'h36 : _GEN_3619; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3621 = 8'h25 == inBytes_14 ? 8'h3f : _GEN_3620; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3622 = 8'h26 == inBytes_14 ? 8'hf7 : _GEN_3621; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3623 = 8'h27 == inBytes_14 ? 8'hcc : _GEN_3622; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3624 = 8'h28 == inBytes_14 ? 8'h34 : _GEN_3623; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3625 = 8'h29 == inBytes_14 ? 8'ha5 : _GEN_3624; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3626 = 8'h2a == inBytes_14 ? 8'he5 : _GEN_3625; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3627 = 8'h2b == inBytes_14 ? 8'hf1 : _GEN_3626; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3628 = 8'h2c == inBytes_14 ? 8'h71 : _GEN_3627; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3629 = 8'h2d == inBytes_14 ? 8'hd8 : _GEN_3628; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3630 = 8'h2e == inBytes_14 ? 8'h31 : _GEN_3629; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3631 = 8'h2f == inBytes_14 ? 8'h15 : _GEN_3630; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3632 = 8'h30 == inBytes_14 ? 8'h4 : _GEN_3631; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3633 = 8'h31 == inBytes_14 ? 8'hc7 : _GEN_3632; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3634 = 8'h32 == inBytes_14 ? 8'h23 : _GEN_3633; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3635 = 8'h33 == inBytes_14 ? 8'hc3 : _GEN_3634; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3636 = 8'h34 == inBytes_14 ? 8'h18 : _GEN_3635; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3637 = 8'h35 == inBytes_14 ? 8'h96 : _GEN_3636; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3638 = 8'h36 == inBytes_14 ? 8'h5 : _GEN_3637; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3639 = 8'h37 == inBytes_14 ? 8'h9a : _GEN_3638; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3640 = 8'h38 == inBytes_14 ? 8'h7 : _GEN_3639; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3641 = 8'h39 == inBytes_14 ? 8'h12 : _GEN_3640; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3642 = 8'h3a == inBytes_14 ? 8'h80 : _GEN_3641; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3643 = 8'h3b == inBytes_14 ? 8'he2 : _GEN_3642; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3644 = 8'h3c == inBytes_14 ? 8'heb : _GEN_3643; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3645 = 8'h3d == inBytes_14 ? 8'h27 : _GEN_3644; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3646 = 8'h3e == inBytes_14 ? 8'hb2 : _GEN_3645; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3647 = 8'h3f == inBytes_14 ? 8'h75 : _GEN_3646; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3648 = 8'h40 == inBytes_14 ? 8'h9 : _GEN_3647; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3649 = 8'h41 == inBytes_14 ? 8'h83 : _GEN_3648; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3650 = 8'h42 == inBytes_14 ? 8'h2c : _GEN_3649; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3651 = 8'h43 == inBytes_14 ? 8'h1a : _GEN_3650; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3652 = 8'h44 == inBytes_14 ? 8'h1b : _GEN_3651; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3653 = 8'h45 == inBytes_14 ? 8'h6e : _GEN_3652; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3654 = 8'h46 == inBytes_14 ? 8'h5a : _GEN_3653; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3655 = 8'h47 == inBytes_14 ? 8'ha0 : _GEN_3654; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3656 = 8'h48 == inBytes_14 ? 8'h52 : _GEN_3655; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3657 = 8'h49 == inBytes_14 ? 8'h3b : _GEN_3656; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3658 = 8'h4a == inBytes_14 ? 8'hd6 : _GEN_3657; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3659 = 8'h4b == inBytes_14 ? 8'hb3 : _GEN_3658; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3660 = 8'h4c == inBytes_14 ? 8'h29 : _GEN_3659; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3661 = 8'h4d == inBytes_14 ? 8'he3 : _GEN_3660; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3662 = 8'h4e == inBytes_14 ? 8'h2f : _GEN_3661; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3663 = 8'h4f == inBytes_14 ? 8'h84 : _GEN_3662; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3664 = 8'h50 == inBytes_14 ? 8'h53 : _GEN_3663; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3665 = 8'h51 == inBytes_14 ? 8'hd1 : _GEN_3664; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3666 = 8'h52 == inBytes_14 ? 8'h0 : _GEN_3665; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3667 = 8'h53 == inBytes_14 ? 8'hed : _GEN_3666; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3668 = 8'h54 == inBytes_14 ? 8'h20 : _GEN_3667; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3669 = 8'h55 == inBytes_14 ? 8'hfc : _GEN_3668; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3670 = 8'h56 == inBytes_14 ? 8'hb1 : _GEN_3669; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3671 = 8'h57 == inBytes_14 ? 8'h5b : _GEN_3670; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3672 = 8'h58 == inBytes_14 ? 8'h6a : _GEN_3671; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3673 = 8'h59 == inBytes_14 ? 8'hcb : _GEN_3672; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3674 = 8'h5a == inBytes_14 ? 8'hbe : _GEN_3673; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3675 = 8'h5b == inBytes_14 ? 8'h39 : _GEN_3674; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3676 = 8'h5c == inBytes_14 ? 8'h4a : _GEN_3675; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3677 = 8'h5d == inBytes_14 ? 8'h4c : _GEN_3676; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3678 = 8'h5e == inBytes_14 ? 8'h58 : _GEN_3677; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3679 = 8'h5f == inBytes_14 ? 8'hcf : _GEN_3678; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3680 = 8'h60 == inBytes_14 ? 8'hd0 : _GEN_3679; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3681 = 8'h61 == inBytes_14 ? 8'hef : _GEN_3680; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3682 = 8'h62 == inBytes_14 ? 8'haa : _GEN_3681; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3683 = 8'h63 == inBytes_14 ? 8'hfb : _GEN_3682; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3684 = 8'h64 == inBytes_14 ? 8'h43 : _GEN_3683; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3685 = 8'h65 == inBytes_14 ? 8'h4d : _GEN_3684; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3686 = 8'h66 == inBytes_14 ? 8'h33 : _GEN_3685; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3687 = 8'h67 == inBytes_14 ? 8'h85 : _GEN_3686; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3688 = 8'h68 == inBytes_14 ? 8'h45 : _GEN_3687; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3689 = 8'h69 == inBytes_14 ? 8'hf9 : _GEN_3688; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3690 = 8'h6a == inBytes_14 ? 8'h2 : _GEN_3689; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3691 = 8'h6b == inBytes_14 ? 8'h7f : _GEN_3690; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3692 = 8'h6c == inBytes_14 ? 8'h50 : _GEN_3691; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3693 = 8'h6d == inBytes_14 ? 8'h3c : _GEN_3692; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3694 = 8'h6e == inBytes_14 ? 8'h9f : _GEN_3693; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3695 = 8'h6f == inBytes_14 ? 8'ha8 : _GEN_3694; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3696 = 8'h70 == inBytes_14 ? 8'h51 : _GEN_3695; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3697 = 8'h71 == inBytes_14 ? 8'ha3 : _GEN_3696; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3698 = 8'h72 == inBytes_14 ? 8'h40 : _GEN_3697; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3699 = 8'h73 == inBytes_14 ? 8'h8f : _GEN_3698; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3700 = 8'h74 == inBytes_14 ? 8'h92 : _GEN_3699; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3701 = 8'h75 == inBytes_14 ? 8'h9d : _GEN_3700; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3702 = 8'h76 == inBytes_14 ? 8'h38 : _GEN_3701; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3703 = 8'h77 == inBytes_14 ? 8'hf5 : _GEN_3702; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3704 = 8'h78 == inBytes_14 ? 8'hbc : _GEN_3703; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3705 = 8'h79 == inBytes_14 ? 8'hb6 : _GEN_3704; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3706 = 8'h7a == inBytes_14 ? 8'hda : _GEN_3705; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3707 = 8'h7b == inBytes_14 ? 8'h21 : _GEN_3706; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3708 = 8'h7c == inBytes_14 ? 8'h10 : _GEN_3707; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3709 = 8'h7d == inBytes_14 ? 8'hff : _GEN_3708; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3710 = 8'h7e == inBytes_14 ? 8'hf3 : _GEN_3709; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3711 = 8'h7f == inBytes_14 ? 8'hd2 : _GEN_3710; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3712 = 8'h80 == inBytes_14 ? 8'hcd : _GEN_3711; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3713 = 8'h81 == inBytes_14 ? 8'hc : _GEN_3712; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3714 = 8'h82 == inBytes_14 ? 8'h13 : _GEN_3713; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3715 = 8'h83 == inBytes_14 ? 8'hec : _GEN_3714; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3716 = 8'h84 == inBytes_14 ? 8'h5f : _GEN_3715; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3717 = 8'h85 == inBytes_14 ? 8'h97 : _GEN_3716; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3718 = 8'h86 == inBytes_14 ? 8'h44 : _GEN_3717; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3719 = 8'h87 == inBytes_14 ? 8'h17 : _GEN_3718; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3720 = 8'h88 == inBytes_14 ? 8'hc4 : _GEN_3719; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3721 = 8'h89 == inBytes_14 ? 8'ha7 : _GEN_3720; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3722 = 8'h8a == inBytes_14 ? 8'h7e : _GEN_3721; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3723 = 8'h8b == inBytes_14 ? 8'h3d : _GEN_3722; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3724 = 8'h8c == inBytes_14 ? 8'h64 : _GEN_3723; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3725 = 8'h8d == inBytes_14 ? 8'h5d : _GEN_3724; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3726 = 8'h8e == inBytes_14 ? 8'h19 : _GEN_3725; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3727 = 8'h8f == inBytes_14 ? 8'h73 : _GEN_3726; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3728 = 8'h90 == inBytes_14 ? 8'h60 : _GEN_3727; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3729 = 8'h91 == inBytes_14 ? 8'h81 : _GEN_3728; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3730 = 8'h92 == inBytes_14 ? 8'h4f : _GEN_3729; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3731 = 8'h93 == inBytes_14 ? 8'hdc : _GEN_3730; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3732 = 8'h94 == inBytes_14 ? 8'h22 : _GEN_3731; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3733 = 8'h95 == inBytes_14 ? 8'h2a : _GEN_3732; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3734 = 8'h96 == inBytes_14 ? 8'h90 : _GEN_3733; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3735 = 8'h97 == inBytes_14 ? 8'h88 : _GEN_3734; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3736 = 8'h98 == inBytes_14 ? 8'h46 : _GEN_3735; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3737 = 8'h99 == inBytes_14 ? 8'hee : _GEN_3736; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3738 = 8'h9a == inBytes_14 ? 8'hb8 : _GEN_3737; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3739 = 8'h9b == inBytes_14 ? 8'h14 : _GEN_3738; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3740 = 8'h9c == inBytes_14 ? 8'hde : _GEN_3739; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3741 = 8'h9d == inBytes_14 ? 8'h5e : _GEN_3740; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3742 = 8'h9e == inBytes_14 ? 8'hb : _GEN_3741; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3743 = 8'h9f == inBytes_14 ? 8'hdb : _GEN_3742; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3744 = 8'ha0 == inBytes_14 ? 8'he0 : _GEN_3743; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3745 = 8'ha1 == inBytes_14 ? 8'h32 : _GEN_3744; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3746 = 8'ha2 == inBytes_14 ? 8'h3a : _GEN_3745; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3747 = 8'ha3 == inBytes_14 ? 8'ha : _GEN_3746; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3748 = 8'ha4 == inBytes_14 ? 8'h49 : _GEN_3747; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3749 = 8'ha5 == inBytes_14 ? 8'h6 : _GEN_3748; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3750 = 8'ha6 == inBytes_14 ? 8'h24 : _GEN_3749; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3751 = 8'ha7 == inBytes_14 ? 8'h5c : _GEN_3750; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3752 = 8'ha8 == inBytes_14 ? 8'hc2 : _GEN_3751; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3753 = 8'ha9 == inBytes_14 ? 8'hd3 : _GEN_3752; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3754 = 8'haa == inBytes_14 ? 8'hac : _GEN_3753; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3755 = 8'hab == inBytes_14 ? 8'h62 : _GEN_3754; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3756 = 8'hac == inBytes_14 ? 8'h91 : _GEN_3755; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3757 = 8'had == inBytes_14 ? 8'h95 : _GEN_3756; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3758 = 8'hae == inBytes_14 ? 8'he4 : _GEN_3757; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3759 = 8'haf == inBytes_14 ? 8'h79 : _GEN_3758; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3760 = 8'hb0 == inBytes_14 ? 8'he7 : _GEN_3759; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3761 = 8'hb1 == inBytes_14 ? 8'hc8 : _GEN_3760; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3762 = 8'hb2 == inBytes_14 ? 8'h37 : _GEN_3761; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3763 = 8'hb3 == inBytes_14 ? 8'h6d : _GEN_3762; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3764 = 8'hb4 == inBytes_14 ? 8'h8d : _GEN_3763; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3765 = 8'hb5 == inBytes_14 ? 8'hd5 : _GEN_3764; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3766 = 8'hb6 == inBytes_14 ? 8'h4e : _GEN_3765; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3767 = 8'hb7 == inBytes_14 ? 8'ha9 : _GEN_3766; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3768 = 8'hb8 == inBytes_14 ? 8'h6c : _GEN_3767; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3769 = 8'hb9 == inBytes_14 ? 8'h56 : _GEN_3768; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3770 = 8'hba == inBytes_14 ? 8'hf4 : _GEN_3769; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3771 = 8'hbb == inBytes_14 ? 8'hea : _GEN_3770; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3772 = 8'hbc == inBytes_14 ? 8'h65 : _GEN_3771; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3773 = 8'hbd == inBytes_14 ? 8'h7a : _GEN_3772; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3774 = 8'hbe == inBytes_14 ? 8'hae : _GEN_3773; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3775 = 8'hbf == inBytes_14 ? 8'h8 : _GEN_3774; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3776 = 8'hc0 == inBytes_14 ? 8'hba : _GEN_3775; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3777 = 8'hc1 == inBytes_14 ? 8'h78 : _GEN_3776; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3778 = 8'hc2 == inBytes_14 ? 8'h25 : _GEN_3777; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3779 = 8'hc3 == inBytes_14 ? 8'h2e : _GEN_3778; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3780 = 8'hc4 == inBytes_14 ? 8'h1c : _GEN_3779; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3781 = 8'hc5 == inBytes_14 ? 8'ha6 : _GEN_3780; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3782 = 8'hc6 == inBytes_14 ? 8'hb4 : _GEN_3781; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3783 = 8'hc7 == inBytes_14 ? 8'hc6 : _GEN_3782; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3784 = 8'hc8 == inBytes_14 ? 8'he8 : _GEN_3783; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3785 = 8'hc9 == inBytes_14 ? 8'hdd : _GEN_3784; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3786 = 8'hca == inBytes_14 ? 8'h74 : _GEN_3785; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3787 = 8'hcb == inBytes_14 ? 8'h1f : _GEN_3786; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3788 = 8'hcc == inBytes_14 ? 8'h4b : _GEN_3787; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3789 = 8'hcd == inBytes_14 ? 8'hbd : _GEN_3788; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3790 = 8'hce == inBytes_14 ? 8'h8b : _GEN_3789; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3791 = 8'hcf == inBytes_14 ? 8'h8a : _GEN_3790; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3792 = 8'hd0 == inBytes_14 ? 8'h70 : _GEN_3791; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3793 = 8'hd1 == inBytes_14 ? 8'h3e : _GEN_3792; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3794 = 8'hd2 == inBytes_14 ? 8'hb5 : _GEN_3793; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3795 = 8'hd3 == inBytes_14 ? 8'h66 : _GEN_3794; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3796 = 8'hd4 == inBytes_14 ? 8'h48 : _GEN_3795; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3797 = 8'hd5 == inBytes_14 ? 8'h3 : _GEN_3796; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3798 = 8'hd6 == inBytes_14 ? 8'hf6 : _GEN_3797; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3799 = 8'hd7 == inBytes_14 ? 8'he : _GEN_3798; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3800 = 8'hd8 == inBytes_14 ? 8'h61 : _GEN_3799; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3801 = 8'hd9 == inBytes_14 ? 8'h35 : _GEN_3800; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3802 = 8'hda == inBytes_14 ? 8'h57 : _GEN_3801; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3803 = 8'hdb == inBytes_14 ? 8'hb9 : _GEN_3802; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3804 = 8'hdc == inBytes_14 ? 8'h86 : _GEN_3803; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3805 = 8'hdd == inBytes_14 ? 8'hc1 : _GEN_3804; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3806 = 8'hde == inBytes_14 ? 8'h1d : _GEN_3805; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3807 = 8'hdf == inBytes_14 ? 8'h9e : _GEN_3806; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3808 = 8'he0 == inBytes_14 ? 8'he1 : _GEN_3807; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3809 = 8'he1 == inBytes_14 ? 8'hf8 : _GEN_3808; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3810 = 8'he2 == inBytes_14 ? 8'h98 : _GEN_3809; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3811 = 8'he3 == inBytes_14 ? 8'h11 : _GEN_3810; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3812 = 8'he4 == inBytes_14 ? 8'h69 : _GEN_3811; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3813 = 8'he5 == inBytes_14 ? 8'hd9 : _GEN_3812; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3814 = 8'he6 == inBytes_14 ? 8'h8e : _GEN_3813; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3815 = 8'he7 == inBytes_14 ? 8'h94 : _GEN_3814; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3816 = 8'he8 == inBytes_14 ? 8'h9b : _GEN_3815; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3817 = 8'he9 == inBytes_14 ? 8'h1e : _GEN_3816; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3818 = 8'hea == inBytes_14 ? 8'h87 : _GEN_3817; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3819 = 8'heb == inBytes_14 ? 8'he9 : _GEN_3818; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3820 = 8'hec == inBytes_14 ? 8'hce : _GEN_3819; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3821 = 8'hed == inBytes_14 ? 8'h55 : _GEN_3820; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3822 = 8'hee == inBytes_14 ? 8'h28 : _GEN_3821; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3823 = 8'hef == inBytes_14 ? 8'hdf : _GEN_3822; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3824 = 8'hf0 == inBytes_14 ? 8'h8c : _GEN_3823; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3825 = 8'hf1 == inBytes_14 ? 8'ha1 : _GEN_3824; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3826 = 8'hf2 == inBytes_14 ? 8'h89 : _GEN_3825; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3827 = 8'hf3 == inBytes_14 ? 8'hd : _GEN_3826; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3828 = 8'hf4 == inBytes_14 ? 8'hbf : _GEN_3827; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3829 = 8'hf5 == inBytes_14 ? 8'he6 : _GEN_3828; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3830 = 8'hf6 == inBytes_14 ? 8'h42 : _GEN_3829; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3831 = 8'hf7 == inBytes_14 ? 8'h68 : _GEN_3830; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3832 = 8'hf8 == inBytes_14 ? 8'h41 : _GEN_3831; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3833 = 8'hf9 == inBytes_14 ? 8'h99 : _GEN_3832; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3834 = 8'hfa == inBytes_14 ? 8'h2d : _GEN_3833; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3835 = 8'hfb == inBytes_14 ? 8'hf : _GEN_3834; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3836 = 8'hfc == inBytes_14 ? 8'hb0 : _GEN_3835; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3837 = 8'hfd == inBytes_14 ? 8'h54 : _GEN_3836; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3838 = 8'hfe == inBytes_14 ? 8'hbb : _GEN_3837; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] outBytes_14 = 8'hff == inBytes_14 ? 8'h16 : _GEN_3838; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3841 = 8'h1 == inBytes_15 ? 8'h7c : 8'h63; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3842 = 8'h2 == inBytes_15 ? 8'h77 : _GEN_3841; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3843 = 8'h3 == inBytes_15 ? 8'h7b : _GEN_3842; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3844 = 8'h4 == inBytes_15 ? 8'hf2 : _GEN_3843; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3845 = 8'h5 == inBytes_15 ? 8'h6b : _GEN_3844; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3846 = 8'h6 == inBytes_15 ? 8'h6f : _GEN_3845; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3847 = 8'h7 == inBytes_15 ? 8'hc5 : _GEN_3846; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3848 = 8'h8 == inBytes_15 ? 8'h30 : _GEN_3847; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3849 = 8'h9 == inBytes_15 ? 8'h1 : _GEN_3848; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3850 = 8'ha == inBytes_15 ? 8'h67 : _GEN_3849; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3851 = 8'hb == inBytes_15 ? 8'h2b : _GEN_3850; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3852 = 8'hc == inBytes_15 ? 8'hfe : _GEN_3851; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3853 = 8'hd == inBytes_15 ? 8'hd7 : _GEN_3852; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3854 = 8'he == inBytes_15 ? 8'hab : _GEN_3853; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3855 = 8'hf == inBytes_15 ? 8'h76 : _GEN_3854; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3856 = 8'h10 == inBytes_15 ? 8'hca : _GEN_3855; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3857 = 8'h11 == inBytes_15 ? 8'h82 : _GEN_3856; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3858 = 8'h12 == inBytes_15 ? 8'hc9 : _GEN_3857; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3859 = 8'h13 == inBytes_15 ? 8'h7d : _GEN_3858; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3860 = 8'h14 == inBytes_15 ? 8'hfa : _GEN_3859; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3861 = 8'h15 == inBytes_15 ? 8'h59 : _GEN_3860; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3862 = 8'h16 == inBytes_15 ? 8'h47 : _GEN_3861; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3863 = 8'h17 == inBytes_15 ? 8'hf0 : _GEN_3862; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3864 = 8'h18 == inBytes_15 ? 8'had : _GEN_3863; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3865 = 8'h19 == inBytes_15 ? 8'hd4 : _GEN_3864; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3866 = 8'h1a == inBytes_15 ? 8'ha2 : _GEN_3865; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3867 = 8'h1b == inBytes_15 ? 8'haf : _GEN_3866; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3868 = 8'h1c == inBytes_15 ? 8'h9c : _GEN_3867; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3869 = 8'h1d == inBytes_15 ? 8'ha4 : _GEN_3868; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3870 = 8'h1e == inBytes_15 ? 8'h72 : _GEN_3869; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3871 = 8'h1f == inBytes_15 ? 8'hc0 : _GEN_3870; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3872 = 8'h20 == inBytes_15 ? 8'hb7 : _GEN_3871; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3873 = 8'h21 == inBytes_15 ? 8'hfd : _GEN_3872; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3874 = 8'h22 == inBytes_15 ? 8'h93 : _GEN_3873; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3875 = 8'h23 == inBytes_15 ? 8'h26 : _GEN_3874; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3876 = 8'h24 == inBytes_15 ? 8'h36 : _GEN_3875; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3877 = 8'h25 == inBytes_15 ? 8'h3f : _GEN_3876; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3878 = 8'h26 == inBytes_15 ? 8'hf7 : _GEN_3877; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3879 = 8'h27 == inBytes_15 ? 8'hcc : _GEN_3878; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3880 = 8'h28 == inBytes_15 ? 8'h34 : _GEN_3879; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3881 = 8'h29 == inBytes_15 ? 8'ha5 : _GEN_3880; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3882 = 8'h2a == inBytes_15 ? 8'he5 : _GEN_3881; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3883 = 8'h2b == inBytes_15 ? 8'hf1 : _GEN_3882; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3884 = 8'h2c == inBytes_15 ? 8'h71 : _GEN_3883; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3885 = 8'h2d == inBytes_15 ? 8'hd8 : _GEN_3884; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3886 = 8'h2e == inBytes_15 ? 8'h31 : _GEN_3885; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3887 = 8'h2f == inBytes_15 ? 8'h15 : _GEN_3886; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3888 = 8'h30 == inBytes_15 ? 8'h4 : _GEN_3887; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3889 = 8'h31 == inBytes_15 ? 8'hc7 : _GEN_3888; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3890 = 8'h32 == inBytes_15 ? 8'h23 : _GEN_3889; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3891 = 8'h33 == inBytes_15 ? 8'hc3 : _GEN_3890; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3892 = 8'h34 == inBytes_15 ? 8'h18 : _GEN_3891; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3893 = 8'h35 == inBytes_15 ? 8'h96 : _GEN_3892; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3894 = 8'h36 == inBytes_15 ? 8'h5 : _GEN_3893; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3895 = 8'h37 == inBytes_15 ? 8'h9a : _GEN_3894; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3896 = 8'h38 == inBytes_15 ? 8'h7 : _GEN_3895; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3897 = 8'h39 == inBytes_15 ? 8'h12 : _GEN_3896; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3898 = 8'h3a == inBytes_15 ? 8'h80 : _GEN_3897; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3899 = 8'h3b == inBytes_15 ? 8'he2 : _GEN_3898; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3900 = 8'h3c == inBytes_15 ? 8'heb : _GEN_3899; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3901 = 8'h3d == inBytes_15 ? 8'h27 : _GEN_3900; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3902 = 8'h3e == inBytes_15 ? 8'hb2 : _GEN_3901; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3903 = 8'h3f == inBytes_15 ? 8'h75 : _GEN_3902; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3904 = 8'h40 == inBytes_15 ? 8'h9 : _GEN_3903; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3905 = 8'h41 == inBytes_15 ? 8'h83 : _GEN_3904; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3906 = 8'h42 == inBytes_15 ? 8'h2c : _GEN_3905; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3907 = 8'h43 == inBytes_15 ? 8'h1a : _GEN_3906; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3908 = 8'h44 == inBytes_15 ? 8'h1b : _GEN_3907; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3909 = 8'h45 == inBytes_15 ? 8'h6e : _GEN_3908; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3910 = 8'h46 == inBytes_15 ? 8'h5a : _GEN_3909; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3911 = 8'h47 == inBytes_15 ? 8'ha0 : _GEN_3910; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3912 = 8'h48 == inBytes_15 ? 8'h52 : _GEN_3911; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3913 = 8'h49 == inBytes_15 ? 8'h3b : _GEN_3912; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3914 = 8'h4a == inBytes_15 ? 8'hd6 : _GEN_3913; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3915 = 8'h4b == inBytes_15 ? 8'hb3 : _GEN_3914; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3916 = 8'h4c == inBytes_15 ? 8'h29 : _GEN_3915; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3917 = 8'h4d == inBytes_15 ? 8'he3 : _GEN_3916; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3918 = 8'h4e == inBytes_15 ? 8'h2f : _GEN_3917; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3919 = 8'h4f == inBytes_15 ? 8'h84 : _GEN_3918; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3920 = 8'h50 == inBytes_15 ? 8'h53 : _GEN_3919; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3921 = 8'h51 == inBytes_15 ? 8'hd1 : _GEN_3920; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3922 = 8'h52 == inBytes_15 ? 8'h0 : _GEN_3921; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3923 = 8'h53 == inBytes_15 ? 8'hed : _GEN_3922; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3924 = 8'h54 == inBytes_15 ? 8'h20 : _GEN_3923; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3925 = 8'h55 == inBytes_15 ? 8'hfc : _GEN_3924; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3926 = 8'h56 == inBytes_15 ? 8'hb1 : _GEN_3925; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3927 = 8'h57 == inBytes_15 ? 8'h5b : _GEN_3926; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3928 = 8'h58 == inBytes_15 ? 8'h6a : _GEN_3927; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3929 = 8'h59 == inBytes_15 ? 8'hcb : _GEN_3928; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3930 = 8'h5a == inBytes_15 ? 8'hbe : _GEN_3929; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3931 = 8'h5b == inBytes_15 ? 8'h39 : _GEN_3930; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3932 = 8'h5c == inBytes_15 ? 8'h4a : _GEN_3931; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3933 = 8'h5d == inBytes_15 ? 8'h4c : _GEN_3932; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3934 = 8'h5e == inBytes_15 ? 8'h58 : _GEN_3933; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3935 = 8'h5f == inBytes_15 ? 8'hcf : _GEN_3934; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3936 = 8'h60 == inBytes_15 ? 8'hd0 : _GEN_3935; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3937 = 8'h61 == inBytes_15 ? 8'hef : _GEN_3936; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3938 = 8'h62 == inBytes_15 ? 8'haa : _GEN_3937; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3939 = 8'h63 == inBytes_15 ? 8'hfb : _GEN_3938; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3940 = 8'h64 == inBytes_15 ? 8'h43 : _GEN_3939; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3941 = 8'h65 == inBytes_15 ? 8'h4d : _GEN_3940; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3942 = 8'h66 == inBytes_15 ? 8'h33 : _GEN_3941; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3943 = 8'h67 == inBytes_15 ? 8'h85 : _GEN_3942; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3944 = 8'h68 == inBytes_15 ? 8'h45 : _GEN_3943; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3945 = 8'h69 == inBytes_15 ? 8'hf9 : _GEN_3944; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3946 = 8'h6a == inBytes_15 ? 8'h2 : _GEN_3945; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3947 = 8'h6b == inBytes_15 ? 8'h7f : _GEN_3946; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3948 = 8'h6c == inBytes_15 ? 8'h50 : _GEN_3947; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3949 = 8'h6d == inBytes_15 ? 8'h3c : _GEN_3948; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3950 = 8'h6e == inBytes_15 ? 8'h9f : _GEN_3949; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3951 = 8'h6f == inBytes_15 ? 8'ha8 : _GEN_3950; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3952 = 8'h70 == inBytes_15 ? 8'h51 : _GEN_3951; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3953 = 8'h71 == inBytes_15 ? 8'ha3 : _GEN_3952; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3954 = 8'h72 == inBytes_15 ? 8'h40 : _GEN_3953; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3955 = 8'h73 == inBytes_15 ? 8'h8f : _GEN_3954; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3956 = 8'h74 == inBytes_15 ? 8'h92 : _GEN_3955; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3957 = 8'h75 == inBytes_15 ? 8'h9d : _GEN_3956; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3958 = 8'h76 == inBytes_15 ? 8'h38 : _GEN_3957; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3959 = 8'h77 == inBytes_15 ? 8'hf5 : _GEN_3958; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3960 = 8'h78 == inBytes_15 ? 8'hbc : _GEN_3959; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3961 = 8'h79 == inBytes_15 ? 8'hb6 : _GEN_3960; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3962 = 8'h7a == inBytes_15 ? 8'hda : _GEN_3961; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3963 = 8'h7b == inBytes_15 ? 8'h21 : _GEN_3962; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3964 = 8'h7c == inBytes_15 ? 8'h10 : _GEN_3963; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3965 = 8'h7d == inBytes_15 ? 8'hff : _GEN_3964; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3966 = 8'h7e == inBytes_15 ? 8'hf3 : _GEN_3965; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3967 = 8'h7f == inBytes_15 ? 8'hd2 : _GEN_3966; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3968 = 8'h80 == inBytes_15 ? 8'hcd : _GEN_3967; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3969 = 8'h81 == inBytes_15 ? 8'hc : _GEN_3968; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3970 = 8'h82 == inBytes_15 ? 8'h13 : _GEN_3969; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3971 = 8'h83 == inBytes_15 ? 8'hec : _GEN_3970; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3972 = 8'h84 == inBytes_15 ? 8'h5f : _GEN_3971; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3973 = 8'h85 == inBytes_15 ? 8'h97 : _GEN_3972; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3974 = 8'h86 == inBytes_15 ? 8'h44 : _GEN_3973; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3975 = 8'h87 == inBytes_15 ? 8'h17 : _GEN_3974; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3976 = 8'h88 == inBytes_15 ? 8'hc4 : _GEN_3975; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3977 = 8'h89 == inBytes_15 ? 8'ha7 : _GEN_3976; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3978 = 8'h8a == inBytes_15 ? 8'h7e : _GEN_3977; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3979 = 8'h8b == inBytes_15 ? 8'h3d : _GEN_3978; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3980 = 8'h8c == inBytes_15 ? 8'h64 : _GEN_3979; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3981 = 8'h8d == inBytes_15 ? 8'h5d : _GEN_3980; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3982 = 8'h8e == inBytes_15 ? 8'h19 : _GEN_3981; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3983 = 8'h8f == inBytes_15 ? 8'h73 : _GEN_3982; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3984 = 8'h90 == inBytes_15 ? 8'h60 : _GEN_3983; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3985 = 8'h91 == inBytes_15 ? 8'h81 : _GEN_3984; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3986 = 8'h92 == inBytes_15 ? 8'h4f : _GEN_3985; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3987 = 8'h93 == inBytes_15 ? 8'hdc : _GEN_3986; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3988 = 8'h94 == inBytes_15 ? 8'h22 : _GEN_3987; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3989 = 8'h95 == inBytes_15 ? 8'h2a : _GEN_3988; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3990 = 8'h96 == inBytes_15 ? 8'h90 : _GEN_3989; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3991 = 8'h97 == inBytes_15 ? 8'h88 : _GEN_3990; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3992 = 8'h98 == inBytes_15 ? 8'h46 : _GEN_3991; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3993 = 8'h99 == inBytes_15 ? 8'hee : _GEN_3992; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3994 = 8'h9a == inBytes_15 ? 8'hb8 : _GEN_3993; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3995 = 8'h9b == inBytes_15 ? 8'h14 : _GEN_3994; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3996 = 8'h9c == inBytes_15 ? 8'hde : _GEN_3995; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3997 = 8'h9d == inBytes_15 ? 8'h5e : _GEN_3996; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3998 = 8'h9e == inBytes_15 ? 8'hb : _GEN_3997; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_3999 = 8'h9f == inBytes_15 ? 8'hdb : _GEN_3998; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_4000 = 8'ha0 == inBytes_15 ? 8'he0 : _GEN_3999; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_4001 = 8'ha1 == inBytes_15 ? 8'h32 : _GEN_4000; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_4002 = 8'ha2 == inBytes_15 ? 8'h3a : _GEN_4001; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_4003 = 8'ha3 == inBytes_15 ? 8'ha : _GEN_4002; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_4004 = 8'ha4 == inBytes_15 ? 8'h49 : _GEN_4003; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_4005 = 8'ha5 == inBytes_15 ? 8'h6 : _GEN_4004; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_4006 = 8'ha6 == inBytes_15 ? 8'h24 : _GEN_4005; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_4007 = 8'ha7 == inBytes_15 ? 8'h5c : _GEN_4006; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_4008 = 8'ha8 == inBytes_15 ? 8'hc2 : _GEN_4007; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_4009 = 8'ha9 == inBytes_15 ? 8'hd3 : _GEN_4008; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_4010 = 8'haa == inBytes_15 ? 8'hac : _GEN_4009; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_4011 = 8'hab == inBytes_15 ? 8'h62 : _GEN_4010; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_4012 = 8'hac == inBytes_15 ? 8'h91 : _GEN_4011; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_4013 = 8'had == inBytes_15 ? 8'h95 : _GEN_4012; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_4014 = 8'hae == inBytes_15 ? 8'he4 : _GEN_4013; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_4015 = 8'haf == inBytes_15 ? 8'h79 : _GEN_4014; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_4016 = 8'hb0 == inBytes_15 ? 8'he7 : _GEN_4015; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_4017 = 8'hb1 == inBytes_15 ? 8'hc8 : _GEN_4016; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_4018 = 8'hb2 == inBytes_15 ? 8'h37 : _GEN_4017; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_4019 = 8'hb3 == inBytes_15 ? 8'h6d : _GEN_4018; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_4020 = 8'hb4 == inBytes_15 ? 8'h8d : _GEN_4019; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_4021 = 8'hb5 == inBytes_15 ? 8'hd5 : _GEN_4020; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_4022 = 8'hb6 == inBytes_15 ? 8'h4e : _GEN_4021; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_4023 = 8'hb7 == inBytes_15 ? 8'ha9 : _GEN_4022; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_4024 = 8'hb8 == inBytes_15 ? 8'h6c : _GEN_4023; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_4025 = 8'hb9 == inBytes_15 ? 8'h56 : _GEN_4024; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_4026 = 8'hba == inBytes_15 ? 8'hf4 : _GEN_4025; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_4027 = 8'hbb == inBytes_15 ? 8'hea : _GEN_4026; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_4028 = 8'hbc == inBytes_15 ? 8'h65 : _GEN_4027; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_4029 = 8'hbd == inBytes_15 ? 8'h7a : _GEN_4028; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_4030 = 8'hbe == inBytes_15 ? 8'hae : _GEN_4029; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_4031 = 8'hbf == inBytes_15 ? 8'h8 : _GEN_4030; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_4032 = 8'hc0 == inBytes_15 ? 8'hba : _GEN_4031; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_4033 = 8'hc1 == inBytes_15 ? 8'h78 : _GEN_4032; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_4034 = 8'hc2 == inBytes_15 ? 8'h25 : _GEN_4033; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_4035 = 8'hc3 == inBytes_15 ? 8'h2e : _GEN_4034; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_4036 = 8'hc4 == inBytes_15 ? 8'h1c : _GEN_4035; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_4037 = 8'hc5 == inBytes_15 ? 8'ha6 : _GEN_4036; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_4038 = 8'hc6 == inBytes_15 ? 8'hb4 : _GEN_4037; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_4039 = 8'hc7 == inBytes_15 ? 8'hc6 : _GEN_4038; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_4040 = 8'hc8 == inBytes_15 ? 8'he8 : _GEN_4039; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_4041 = 8'hc9 == inBytes_15 ? 8'hdd : _GEN_4040; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_4042 = 8'hca == inBytes_15 ? 8'h74 : _GEN_4041; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_4043 = 8'hcb == inBytes_15 ? 8'h1f : _GEN_4042; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_4044 = 8'hcc == inBytes_15 ? 8'h4b : _GEN_4043; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_4045 = 8'hcd == inBytes_15 ? 8'hbd : _GEN_4044; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_4046 = 8'hce == inBytes_15 ? 8'h8b : _GEN_4045; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_4047 = 8'hcf == inBytes_15 ? 8'h8a : _GEN_4046; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_4048 = 8'hd0 == inBytes_15 ? 8'h70 : _GEN_4047; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_4049 = 8'hd1 == inBytes_15 ? 8'h3e : _GEN_4048; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_4050 = 8'hd2 == inBytes_15 ? 8'hb5 : _GEN_4049; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_4051 = 8'hd3 == inBytes_15 ? 8'h66 : _GEN_4050; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_4052 = 8'hd4 == inBytes_15 ? 8'h48 : _GEN_4051; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_4053 = 8'hd5 == inBytes_15 ? 8'h3 : _GEN_4052; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_4054 = 8'hd6 == inBytes_15 ? 8'hf6 : _GEN_4053; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_4055 = 8'hd7 == inBytes_15 ? 8'he : _GEN_4054; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_4056 = 8'hd8 == inBytes_15 ? 8'h61 : _GEN_4055; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_4057 = 8'hd9 == inBytes_15 ? 8'h35 : _GEN_4056; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_4058 = 8'hda == inBytes_15 ? 8'h57 : _GEN_4057; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_4059 = 8'hdb == inBytes_15 ? 8'hb9 : _GEN_4058; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_4060 = 8'hdc == inBytes_15 ? 8'h86 : _GEN_4059; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_4061 = 8'hdd == inBytes_15 ? 8'hc1 : _GEN_4060; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_4062 = 8'hde == inBytes_15 ? 8'h1d : _GEN_4061; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_4063 = 8'hdf == inBytes_15 ? 8'h9e : _GEN_4062; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_4064 = 8'he0 == inBytes_15 ? 8'he1 : _GEN_4063; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_4065 = 8'he1 == inBytes_15 ? 8'hf8 : _GEN_4064; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_4066 = 8'he2 == inBytes_15 ? 8'h98 : _GEN_4065; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_4067 = 8'he3 == inBytes_15 ? 8'h11 : _GEN_4066; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_4068 = 8'he4 == inBytes_15 ? 8'h69 : _GEN_4067; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_4069 = 8'he5 == inBytes_15 ? 8'hd9 : _GEN_4068; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_4070 = 8'he6 == inBytes_15 ? 8'h8e : _GEN_4069; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_4071 = 8'he7 == inBytes_15 ? 8'h94 : _GEN_4070; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_4072 = 8'he8 == inBytes_15 ? 8'h9b : _GEN_4071; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_4073 = 8'he9 == inBytes_15 ? 8'h1e : _GEN_4072; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_4074 = 8'hea == inBytes_15 ? 8'h87 : _GEN_4073; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_4075 = 8'heb == inBytes_15 ? 8'he9 : _GEN_4074; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_4076 = 8'hec == inBytes_15 ? 8'hce : _GEN_4075; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_4077 = 8'hed == inBytes_15 ? 8'h55 : _GEN_4076; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_4078 = 8'hee == inBytes_15 ? 8'h28 : _GEN_4077; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_4079 = 8'hef == inBytes_15 ? 8'hdf : _GEN_4078; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_4080 = 8'hf0 == inBytes_15 ? 8'h8c : _GEN_4079; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_4081 = 8'hf1 == inBytes_15 ? 8'ha1 : _GEN_4080; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_4082 = 8'hf2 == inBytes_15 ? 8'h89 : _GEN_4081; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_4083 = 8'hf3 == inBytes_15 ? 8'hd : _GEN_4082; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_4084 = 8'hf4 == inBytes_15 ? 8'hbf : _GEN_4083; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_4085 = 8'hf5 == inBytes_15 ? 8'he6 : _GEN_4084; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_4086 = 8'hf6 == inBytes_15 ? 8'h42 : _GEN_4085; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_4087 = 8'hf7 == inBytes_15 ? 8'h68 : _GEN_4086; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_4088 = 8'hf8 == inBytes_15 ? 8'h41 : _GEN_4087; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_4089 = 8'hf9 == inBytes_15 ? 8'h99 : _GEN_4088; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_4090 = 8'hfa == inBytes_15 ? 8'h2d : _GEN_4089; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_4091 = 8'hfb == inBytes_15 ? 8'hf : _GEN_4090; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_4092 = 8'hfc == inBytes_15 ? 8'hb0 : _GEN_4091; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_4093 = 8'hfd == inBytes_15 ? 8'h54 : _GEN_4092; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] _GEN_4094 = 8'hfe == inBytes_15 ? 8'hbb : _GEN_4093; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [7:0] outBytes_15 = 8'hff == inBytes_15 ? 8'h16 : _GEN_4094; // @[src/main/scala/crypto/aes/SubBytes.scala 58:{39,39}]
  wire [63:0] outWord_lo = {outBytes_8,outBytes_9,outBytes_10,outBytes_11,outBytes_12,outBytes_13,outBytes_14,
    outBytes_15}; // @[src/main/scala/crypto/aes/SubBytes.scala 60:20]
  wire [63:0] outWord_hi = {outBytes_0,outBytes_1,outBytes_2,outBytes_3,outBytes_4,outBytes_5,outBytes_6,outBytes_7}; // @[src/main/scala/crypto/aes/SubBytes.scala 60:20]
  assign io_in_ready = io_out_ready; // @[src/main/scala/crypto/aes/SubBytes.scala 15:16]
  assign io_out_valid = io_in_valid; // @[src/main/scala/crypto/aes/SubBytes.scala 14:16]
  assign io_out_bits_bits = {outWord_hi,outWord_lo}; // @[src/main/scala/crypto/aes/SubBytes.scala 60:20]
endmodule
module ShiftRows(
  output         io_in_ready, // @[src/main/scala/crypto/aes/ShiftRows.scala 9:14]
  input          io_in_valid, // @[src/main/scala/crypto/aes/ShiftRows.scala 9:14]
  input  [127:0] io_in_bits_bits, // @[src/main/scala/crypto/aes/ShiftRows.scala 9:14]
  input          io_out_ready, // @[src/main/scala/crypto/aes/ShiftRows.scala 9:14]
  output         io_out_valid, // @[src/main/scala/crypto/aes/ShiftRows.scala 9:14]
  output [127:0] io_out_bits_bits // @[src/main/scala/crypto/aes/ShiftRows.scala 9:14]
);
  wire [7:0] bytes_0 = io_in_bits_bits[127:120]; // @[src/main/scala/crypto/aes/ShiftRows.scala 21:39]
  wire [7:0] bytes_1 = io_in_bits_bits[119:112]; // @[src/main/scala/crypto/aes/ShiftRows.scala 21:39]
  wire [7:0] bytes_2 = io_in_bits_bits[111:104]; // @[src/main/scala/crypto/aes/ShiftRows.scala 21:39]
  wire [7:0] bytes_3 = io_in_bits_bits[103:96]; // @[src/main/scala/crypto/aes/ShiftRows.scala 21:39]
  wire [7:0] bytes_4 = io_in_bits_bits[95:88]; // @[src/main/scala/crypto/aes/ShiftRows.scala 21:39]
  wire [7:0] bytes_5 = io_in_bits_bits[87:80]; // @[src/main/scala/crypto/aes/ShiftRows.scala 21:39]
  wire [7:0] bytes_6 = io_in_bits_bits[79:72]; // @[src/main/scala/crypto/aes/ShiftRows.scala 21:39]
  wire [7:0] bytes_7 = io_in_bits_bits[71:64]; // @[src/main/scala/crypto/aes/ShiftRows.scala 21:39]
  wire [7:0] bytes_8 = io_in_bits_bits[63:56]; // @[src/main/scala/crypto/aes/ShiftRows.scala 21:39]
  wire [7:0] bytes_9 = io_in_bits_bits[55:48]; // @[src/main/scala/crypto/aes/ShiftRows.scala 21:39]
  wire [7:0] bytes_10 = io_in_bits_bits[47:40]; // @[src/main/scala/crypto/aes/ShiftRows.scala 21:39]
  wire [7:0] bytes_11 = io_in_bits_bits[39:32]; // @[src/main/scala/crypto/aes/ShiftRows.scala 21:39]
  wire [7:0] bytes_12 = io_in_bits_bits[31:24]; // @[src/main/scala/crypto/aes/ShiftRows.scala 21:39]
  wire [7:0] bytes_13 = io_in_bits_bits[23:16]; // @[src/main/scala/crypto/aes/ShiftRows.scala 21:39]
  wire [7:0] bytes_14 = io_in_bits_bits[15:8]; // @[src/main/scala/crypto/aes/ShiftRows.scala 21:39]
  wire [7:0] bytes_15 = io_in_bits_bits[7:0]; // @[src/main/scala/crypto/aes/ShiftRows.scala 21:39]
  wire [63:0] outWord_lo = {bytes_8,bytes_13,bytes_2,bytes_7,bytes_12,bytes_1,bytes_6,bytes_11}; // @[src/main/scala/crypto/aes/ShiftRows.scala 48:20]
  wire [63:0] outWord_hi = {bytes_0,bytes_5,bytes_10,bytes_15,bytes_4,bytes_9,bytes_14,bytes_3}; // @[src/main/scala/crypto/aes/ShiftRows.scala 48:20]
  assign io_in_ready = io_out_ready; // @[src/main/scala/crypto/aes/ShiftRows.scala 16:16]
  assign io_out_valid = io_in_valid; // @[src/main/scala/crypto/aes/ShiftRows.scala 15:16]
  assign io_out_bits_bits = {outWord_hi,outWord_lo}; // @[src/main/scala/crypto/aes/ShiftRows.scala 48:20]
endmodule
module MixColumns(
  output         io_in_ready, // @[src/main/scala/crypto/aes/MixColumns.scala 9:14]
  input          io_in_valid, // @[src/main/scala/crypto/aes/MixColumns.scala 9:14]
  input  [127:0] io_in_bits_bits, // @[src/main/scala/crypto/aes/MixColumns.scala 9:14]
  input          io_out_ready, // @[src/main/scala/crypto/aes/MixColumns.scala 9:14]
  output         io_out_valid, // @[src/main/scala/crypto/aes/MixColumns.scala 9:14]
  output [127:0] io_out_bits_bits // @[src/main/scala/crypto/aes/MixColumns.scala 9:14]
);
  wire [7:0] bytes_0 = io_in_bits_bits[127:120]; // @[src/main/scala/crypto/aes/MixColumns.scala 19:40]
  wire [7:0] bytes_1 = io_in_bits_bits[119:112]; // @[src/main/scala/crypto/aes/MixColumns.scala 19:40]
  wire [7:0] bytes_2 = io_in_bits_bits[111:104]; // @[src/main/scala/crypto/aes/MixColumns.scala 19:40]
  wire [7:0] bytes_3 = io_in_bits_bits[103:96]; // @[src/main/scala/crypto/aes/MixColumns.scala 19:40]
  wire [7:0] bytes_4 = io_in_bits_bits[95:88]; // @[src/main/scala/crypto/aes/MixColumns.scala 19:40]
  wire [7:0] bytes_5 = io_in_bits_bits[87:80]; // @[src/main/scala/crypto/aes/MixColumns.scala 19:40]
  wire [7:0] bytes_6 = io_in_bits_bits[79:72]; // @[src/main/scala/crypto/aes/MixColumns.scala 19:40]
  wire [7:0] bytes_7 = io_in_bits_bits[71:64]; // @[src/main/scala/crypto/aes/MixColumns.scala 19:40]
  wire [7:0] bytes_8 = io_in_bits_bits[63:56]; // @[src/main/scala/crypto/aes/MixColumns.scala 19:40]
  wire [7:0] bytes_9 = io_in_bits_bits[55:48]; // @[src/main/scala/crypto/aes/MixColumns.scala 19:40]
  wire [7:0] bytes_10 = io_in_bits_bits[47:40]; // @[src/main/scala/crypto/aes/MixColumns.scala 19:40]
  wire [7:0] bytes_11 = io_in_bits_bits[39:32]; // @[src/main/scala/crypto/aes/MixColumns.scala 19:40]
  wire [7:0] bytes_12 = io_in_bits_bits[31:24]; // @[src/main/scala/crypto/aes/MixColumns.scala 19:40]
  wire [7:0] bytes_13 = io_in_bits_bits[23:16]; // @[src/main/scala/crypto/aes/MixColumns.scala 19:40]
  wire [7:0] bytes_14 = io_in_bits_bits[15:8]; // @[src/main/scala/crypto/aes/MixColumns.scala 19:40]
  wire [7:0] bytes_15 = io_in_bits_bits[7:0]; // @[src/main/scala/crypto/aes/MixColumns.scala 19:40]
  wire  r0_msb = bytes_0[7]; // @[src/main/scala/crypto/aes/MixColumns.scala 22:16]
  wire [8:0] _r0_sh_T = {bytes_0, 1'h0}; // @[src/main/scala/crypto/aes/MixColumns.scala 23:18]
  wire [7:0] r0_sh = _r0_sh_T[7:0]; // @[src/main/scala/crypto/aes/MixColumns.scala 23:23]
  wire [7:0] _r0_T = r0_sh ^ 8'h1b; // @[src/main/scala/crypto/aes/MixColumns.scala 24:17]
  wire [7:0] _r0_T_1 = r0_msb ? _r0_T : r0_sh; // @[src/main/scala/crypto/aes/MixColumns.scala 24:8]
  wire  r0_msb_1 = bytes_1[7]; // @[src/main/scala/crypto/aes/MixColumns.scala 22:16]
  wire [8:0] _r0_sh_T_1 = {bytes_1, 1'h0}; // @[src/main/scala/crypto/aes/MixColumns.scala 23:18]
  wire [7:0] r0_sh_1 = _r0_sh_T_1[7:0]; // @[src/main/scala/crypto/aes/MixColumns.scala 23:23]
  wire [7:0] _r0_T_2 = r0_sh_1 ^ 8'h1b; // @[src/main/scala/crypto/aes/MixColumns.scala 24:17]
  wire [7:0] _r0_T_3 = r0_msb_1 ? _r0_T_2 : r0_sh_1; // @[src/main/scala/crypto/aes/MixColumns.scala 24:8]
  wire [7:0] _r0_T_4 = _r0_T_3 ^ bytes_1; // @[src/main/scala/crypto/aes/MixColumns.scala 27:38]
  wire [7:0] _r0_T_5 = _r0_T_1 ^ _r0_T_4; // @[src/main/scala/crypto/aes/MixColumns.scala 31:23]
  wire [7:0] _r0_T_6 = _r0_T_5 ^ bytes_2; // @[src/main/scala/crypto/aes/MixColumns.scala 31:34]
  wire [7:0] r0 = _r0_T_6 ^ bytes_3; // @[src/main/scala/crypto/aes/MixColumns.scala 31:45]
  wire [7:0] _r1_T_2 = bytes_0 ^ _r0_T_3; // @[src/main/scala/crypto/aes/MixColumns.scala 32:23]
  wire  r1_msb_1 = bytes_2[7]; // @[src/main/scala/crypto/aes/MixColumns.scala 22:16]
  wire [8:0] _r1_sh_T_1 = {bytes_2, 1'h0}; // @[src/main/scala/crypto/aes/MixColumns.scala 23:18]
  wire [7:0] r1_sh_1 = _r1_sh_T_1[7:0]; // @[src/main/scala/crypto/aes/MixColumns.scala 23:23]
  wire [7:0] _r1_T_3 = r1_sh_1 ^ 8'h1b; // @[src/main/scala/crypto/aes/MixColumns.scala 24:17]
  wire [7:0] _r1_T_4 = r1_msb_1 ? _r1_T_3 : r1_sh_1; // @[src/main/scala/crypto/aes/MixColumns.scala 24:8]
  wire [7:0] _r1_T_5 = _r1_T_4 ^ bytes_2; // @[src/main/scala/crypto/aes/MixColumns.scala 27:38]
  wire [7:0] _r1_T_6 = _r1_T_2 ^ _r1_T_5; // @[src/main/scala/crypto/aes/MixColumns.scala 32:34]
  wire [7:0] r1 = _r1_T_6 ^ bytes_3; // @[src/main/scala/crypto/aes/MixColumns.scala 32:45]
  wire [7:0] _r2_T = bytes_0 ^ bytes_1; // @[src/main/scala/crypto/aes/MixColumns.scala 33:23]
  wire [7:0] _r2_T_3 = _r2_T ^ _r1_T_4; // @[src/main/scala/crypto/aes/MixColumns.scala 33:34]
  wire  r2_msb_1 = bytes_3[7]; // @[src/main/scala/crypto/aes/MixColumns.scala 22:16]
  wire [8:0] _r2_sh_T_1 = {bytes_3, 1'h0}; // @[src/main/scala/crypto/aes/MixColumns.scala 23:18]
  wire [7:0] r2_sh_1 = _r2_sh_T_1[7:0]; // @[src/main/scala/crypto/aes/MixColumns.scala 23:23]
  wire [7:0] _r2_T_4 = r2_sh_1 ^ 8'h1b; // @[src/main/scala/crypto/aes/MixColumns.scala 24:17]
  wire [7:0] _r2_T_5 = r2_msb_1 ? _r2_T_4 : r2_sh_1; // @[src/main/scala/crypto/aes/MixColumns.scala 24:8]
  wire [7:0] _r2_T_6 = _r2_T_5 ^ bytes_3; // @[src/main/scala/crypto/aes/MixColumns.scala 27:38]
  wire [7:0] r2 = _r2_T_3 ^ _r2_T_6; // @[src/main/scala/crypto/aes/MixColumns.scala 33:45]
  wire [7:0] _r3_T_2 = _r0_T_1 ^ bytes_0; // @[src/main/scala/crypto/aes/MixColumns.scala 27:38]
  wire [7:0] _r3_T_3 = _r3_T_2 ^ bytes_1; // @[src/main/scala/crypto/aes/MixColumns.scala 34:23]
  wire [7:0] _r3_T_4 = _r3_T_3 ^ bytes_2; // @[src/main/scala/crypto/aes/MixColumns.scala 34:34]
  wire [7:0] r3 = _r3_T_4 ^ _r2_T_5; // @[src/main/scala/crypto/aes/MixColumns.scala 34:45]
  wire  r0_msb_2 = bytes_4[7]; // @[src/main/scala/crypto/aes/MixColumns.scala 22:16]
  wire [8:0] _r0_sh_T_2 = {bytes_4, 1'h0}; // @[src/main/scala/crypto/aes/MixColumns.scala 23:18]
  wire [7:0] r0_sh_2 = _r0_sh_T_2[7:0]; // @[src/main/scala/crypto/aes/MixColumns.scala 23:23]
  wire [7:0] _r0_T_7 = r0_sh_2 ^ 8'h1b; // @[src/main/scala/crypto/aes/MixColumns.scala 24:17]
  wire [7:0] _r0_T_8 = r0_msb_2 ? _r0_T_7 : r0_sh_2; // @[src/main/scala/crypto/aes/MixColumns.scala 24:8]
  wire  r0_msb_3 = bytes_5[7]; // @[src/main/scala/crypto/aes/MixColumns.scala 22:16]
  wire [8:0] _r0_sh_T_3 = {bytes_5, 1'h0}; // @[src/main/scala/crypto/aes/MixColumns.scala 23:18]
  wire [7:0] r0_sh_3 = _r0_sh_T_3[7:0]; // @[src/main/scala/crypto/aes/MixColumns.scala 23:23]
  wire [7:0] _r0_T_9 = r0_sh_3 ^ 8'h1b; // @[src/main/scala/crypto/aes/MixColumns.scala 24:17]
  wire [7:0] _r0_T_10 = r0_msb_3 ? _r0_T_9 : r0_sh_3; // @[src/main/scala/crypto/aes/MixColumns.scala 24:8]
  wire [7:0] _r0_T_11 = _r0_T_10 ^ bytes_5; // @[src/main/scala/crypto/aes/MixColumns.scala 27:38]
  wire [7:0] _r0_T_12 = _r0_T_8 ^ _r0_T_11; // @[src/main/scala/crypto/aes/MixColumns.scala 31:23]
  wire [7:0] _r0_T_13 = _r0_T_12 ^ bytes_6; // @[src/main/scala/crypto/aes/MixColumns.scala 31:34]
  wire [7:0] r0_1 = _r0_T_13 ^ bytes_7; // @[src/main/scala/crypto/aes/MixColumns.scala 31:45]
  wire [7:0] _r1_T_9 = bytes_4 ^ _r0_T_10; // @[src/main/scala/crypto/aes/MixColumns.scala 32:23]
  wire  r1_msb_3 = bytes_6[7]; // @[src/main/scala/crypto/aes/MixColumns.scala 22:16]
  wire [8:0] _r1_sh_T_3 = {bytes_6, 1'h0}; // @[src/main/scala/crypto/aes/MixColumns.scala 23:18]
  wire [7:0] r1_sh_3 = _r1_sh_T_3[7:0]; // @[src/main/scala/crypto/aes/MixColumns.scala 23:23]
  wire [7:0] _r1_T_10 = r1_sh_3 ^ 8'h1b; // @[src/main/scala/crypto/aes/MixColumns.scala 24:17]
  wire [7:0] _r1_T_11 = r1_msb_3 ? _r1_T_10 : r1_sh_3; // @[src/main/scala/crypto/aes/MixColumns.scala 24:8]
  wire [7:0] _r1_T_12 = _r1_T_11 ^ bytes_6; // @[src/main/scala/crypto/aes/MixColumns.scala 27:38]
  wire [7:0] _r1_T_13 = _r1_T_9 ^ _r1_T_12; // @[src/main/scala/crypto/aes/MixColumns.scala 32:34]
  wire [7:0] r1_1 = _r1_T_13 ^ bytes_7; // @[src/main/scala/crypto/aes/MixColumns.scala 32:45]
  wire [7:0] _r2_T_7 = bytes_4 ^ bytes_5; // @[src/main/scala/crypto/aes/MixColumns.scala 33:23]
  wire [7:0] _r2_T_10 = _r2_T_7 ^ _r1_T_11; // @[src/main/scala/crypto/aes/MixColumns.scala 33:34]
  wire  r2_msb_3 = bytes_7[7]; // @[src/main/scala/crypto/aes/MixColumns.scala 22:16]
  wire [8:0] _r2_sh_T_3 = {bytes_7, 1'h0}; // @[src/main/scala/crypto/aes/MixColumns.scala 23:18]
  wire [7:0] r2_sh_3 = _r2_sh_T_3[7:0]; // @[src/main/scala/crypto/aes/MixColumns.scala 23:23]
  wire [7:0] _r2_T_11 = r2_sh_3 ^ 8'h1b; // @[src/main/scala/crypto/aes/MixColumns.scala 24:17]
  wire [7:0] _r2_T_12 = r2_msb_3 ? _r2_T_11 : r2_sh_3; // @[src/main/scala/crypto/aes/MixColumns.scala 24:8]
  wire [7:0] _r2_T_13 = _r2_T_12 ^ bytes_7; // @[src/main/scala/crypto/aes/MixColumns.scala 27:38]
  wire [7:0] r2_1 = _r2_T_10 ^ _r2_T_13; // @[src/main/scala/crypto/aes/MixColumns.scala 33:45]
  wire [7:0] _r3_T_9 = _r0_T_8 ^ bytes_4; // @[src/main/scala/crypto/aes/MixColumns.scala 27:38]
  wire [7:0] _r3_T_10 = _r3_T_9 ^ bytes_5; // @[src/main/scala/crypto/aes/MixColumns.scala 34:23]
  wire [7:0] _r3_T_11 = _r3_T_10 ^ bytes_6; // @[src/main/scala/crypto/aes/MixColumns.scala 34:34]
  wire [7:0] r3_1 = _r3_T_11 ^ _r2_T_12; // @[src/main/scala/crypto/aes/MixColumns.scala 34:45]
  wire  r0_msb_4 = bytes_8[7]; // @[src/main/scala/crypto/aes/MixColumns.scala 22:16]
  wire [8:0] _r0_sh_T_4 = {bytes_8, 1'h0}; // @[src/main/scala/crypto/aes/MixColumns.scala 23:18]
  wire [7:0] r0_sh_4 = _r0_sh_T_4[7:0]; // @[src/main/scala/crypto/aes/MixColumns.scala 23:23]
  wire [7:0] _r0_T_14 = r0_sh_4 ^ 8'h1b; // @[src/main/scala/crypto/aes/MixColumns.scala 24:17]
  wire [7:0] _r0_T_15 = r0_msb_4 ? _r0_T_14 : r0_sh_4; // @[src/main/scala/crypto/aes/MixColumns.scala 24:8]
  wire  r0_msb_5 = bytes_9[7]; // @[src/main/scala/crypto/aes/MixColumns.scala 22:16]
  wire [8:0] _r0_sh_T_5 = {bytes_9, 1'h0}; // @[src/main/scala/crypto/aes/MixColumns.scala 23:18]
  wire [7:0] r0_sh_5 = _r0_sh_T_5[7:0]; // @[src/main/scala/crypto/aes/MixColumns.scala 23:23]
  wire [7:0] _r0_T_16 = r0_sh_5 ^ 8'h1b; // @[src/main/scala/crypto/aes/MixColumns.scala 24:17]
  wire [7:0] _r0_T_17 = r0_msb_5 ? _r0_T_16 : r0_sh_5; // @[src/main/scala/crypto/aes/MixColumns.scala 24:8]
  wire [7:0] _r0_T_18 = _r0_T_17 ^ bytes_9; // @[src/main/scala/crypto/aes/MixColumns.scala 27:38]
  wire [7:0] _r0_T_19 = _r0_T_15 ^ _r0_T_18; // @[src/main/scala/crypto/aes/MixColumns.scala 31:23]
  wire [7:0] _r0_T_20 = _r0_T_19 ^ bytes_10; // @[src/main/scala/crypto/aes/MixColumns.scala 31:34]
  wire [7:0] r0_2 = _r0_T_20 ^ bytes_11; // @[src/main/scala/crypto/aes/MixColumns.scala 31:45]
  wire [7:0] _r1_T_16 = bytes_8 ^ _r0_T_17; // @[src/main/scala/crypto/aes/MixColumns.scala 32:23]
  wire  r1_msb_5 = bytes_10[7]; // @[src/main/scala/crypto/aes/MixColumns.scala 22:16]
  wire [8:0] _r1_sh_T_5 = {bytes_10, 1'h0}; // @[src/main/scala/crypto/aes/MixColumns.scala 23:18]
  wire [7:0] r1_sh_5 = _r1_sh_T_5[7:0]; // @[src/main/scala/crypto/aes/MixColumns.scala 23:23]
  wire [7:0] _r1_T_17 = r1_sh_5 ^ 8'h1b; // @[src/main/scala/crypto/aes/MixColumns.scala 24:17]
  wire [7:0] _r1_T_18 = r1_msb_5 ? _r1_T_17 : r1_sh_5; // @[src/main/scala/crypto/aes/MixColumns.scala 24:8]
  wire [7:0] _r1_T_19 = _r1_T_18 ^ bytes_10; // @[src/main/scala/crypto/aes/MixColumns.scala 27:38]
  wire [7:0] _r1_T_20 = _r1_T_16 ^ _r1_T_19; // @[src/main/scala/crypto/aes/MixColumns.scala 32:34]
  wire [7:0] r1_2 = _r1_T_20 ^ bytes_11; // @[src/main/scala/crypto/aes/MixColumns.scala 32:45]
  wire [7:0] _r2_T_14 = bytes_8 ^ bytes_9; // @[src/main/scala/crypto/aes/MixColumns.scala 33:23]
  wire [7:0] _r2_T_17 = _r2_T_14 ^ _r1_T_18; // @[src/main/scala/crypto/aes/MixColumns.scala 33:34]
  wire  r2_msb_5 = bytes_11[7]; // @[src/main/scala/crypto/aes/MixColumns.scala 22:16]
  wire [8:0] _r2_sh_T_5 = {bytes_11, 1'h0}; // @[src/main/scala/crypto/aes/MixColumns.scala 23:18]
  wire [7:0] r2_sh_5 = _r2_sh_T_5[7:0]; // @[src/main/scala/crypto/aes/MixColumns.scala 23:23]
  wire [7:0] _r2_T_18 = r2_sh_5 ^ 8'h1b; // @[src/main/scala/crypto/aes/MixColumns.scala 24:17]
  wire [7:0] _r2_T_19 = r2_msb_5 ? _r2_T_18 : r2_sh_5; // @[src/main/scala/crypto/aes/MixColumns.scala 24:8]
  wire [7:0] _r2_T_20 = _r2_T_19 ^ bytes_11; // @[src/main/scala/crypto/aes/MixColumns.scala 27:38]
  wire [7:0] r2_2 = _r2_T_17 ^ _r2_T_20; // @[src/main/scala/crypto/aes/MixColumns.scala 33:45]
  wire [7:0] _r3_T_16 = _r0_T_15 ^ bytes_8; // @[src/main/scala/crypto/aes/MixColumns.scala 27:38]
  wire [7:0] _r3_T_17 = _r3_T_16 ^ bytes_9; // @[src/main/scala/crypto/aes/MixColumns.scala 34:23]
  wire [7:0] _r3_T_18 = _r3_T_17 ^ bytes_10; // @[src/main/scala/crypto/aes/MixColumns.scala 34:34]
  wire [7:0] r3_2 = _r3_T_18 ^ _r2_T_19; // @[src/main/scala/crypto/aes/MixColumns.scala 34:45]
  wire  r0_msb_6 = bytes_12[7]; // @[src/main/scala/crypto/aes/MixColumns.scala 22:16]
  wire [8:0] _r0_sh_T_6 = {bytes_12, 1'h0}; // @[src/main/scala/crypto/aes/MixColumns.scala 23:18]
  wire [7:0] r0_sh_6 = _r0_sh_T_6[7:0]; // @[src/main/scala/crypto/aes/MixColumns.scala 23:23]
  wire [7:0] _r0_T_21 = r0_sh_6 ^ 8'h1b; // @[src/main/scala/crypto/aes/MixColumns.scala 24:17]
  wire [7:0] _r0_T_22 = r0_msb_6 ? _r0_T_21 : r0_sh_6; // @[src/main/scala/crypto/aes/MixColumns.scala 24:8]
  wire  r0_msb_7 = bytes_13[7]; // @[src/main/scala/crypto/aes/MixColumns.scala 22:16]
  wire [8:0] _r0_sh_T_7 = {bytes_13, 1'h0}; // @[src/main/scala/crypto/aes/MixColumns.scala 23:18]
  wire [7:0] r0_sh_7 = _r0_sh_T_7[7:0]; // @[src/main/scala/crypto/aes/MixColumns.scala 23:23]
  wire [7:0] _r0_T_23 = r0_sh_7 ^ 8'h1b; // @[src/main/scala/crypto/aes/MixColumns.scala 24:17]
  wire [7:0] _r0_T_24 = r0_msb_7 ? _r0_T_23 : r0_sh_7; // @[src/main/scala/crypto/aes/MixColumns.scala 24:8]
  wire [7:0] _r0_T_25 = _r0_T_24 ^ bytes_13; // @[src/main/scala/crypto/aes/MixColumns.scala 27:38]
  wire [7:0] _r0_T_26 = _r0_T_22 ^ _r0_T_25; // @[src/main/scala/crypto/aes/MixColumns.scala 31:23]
  wire [7:0] _r0_T_27 = _r0_T_26 ^ bytes_14; // @[src/main/scala/crypto/aes/MixColumns.scala 31:34]
  wire [7:0] r0_3 = _r0_T_27 ^ bytes_15; // @[src/main/scala/crypto/aes/MixColumns.scala 31:45]
  wire [7:0] _r1_T_23 = bytes_12 ^ _r0_T_24; // @[src/main/scala/crypto/aes/MixColumns.scala 32:23]
  wire  r1_msb_7 = bytes_14[7]; // @[src/main/scala/crypto/aes/MixColumns.scala 22:16]
  wire [8:0] _r1_sh_T_7 = {bytes_14, 1'h0}; // @[src/main/scala/crypto/aes/MixColumns.scala 23:18]
  wire [7:0] r1_sh_7 = _r1_sh_T_7[7:0]; // @[src/main/scala/crypto/aes/MixColumns.scala 23:23]
  wire [7:0] _r1_T_24 = r1_sh_7 ^ 8'h1b; // @[src/main/scala/crypto/aes/MixColumns.scala 24:17]
  wire [7:0] _r1_T_25 = r1_msb_7 ? _r1_T_24 : r1_sh_7; // @[src/main/scala/crypto/aes/MixColumns.scala 24:8]
  wire [7:0] _r1_T_26 = _r1_T_25 ^ bytes_14; // @[src/main/scala/crypto/aes/MixColumns.scala 27:38]
  wire [7:0] _r1_T_27 = _r1_T_23 ^ _r1_T_26; // @[src/main/scala/crypto/aes/MixColumns.scala 32:34]
  wire [7:0] r1_3 = _r1_T_27 ^ bytes_15; // @[src/main/scala/crypto/aes/MixColumns.scala 32:45]
  wire [7:0] _r2_T_21 = bytes_12 ^ bytes_13; // @[src/main/scala/crypto/aes/MixColumns.scala 33:23]
  wire [7:0] _r2_T_24 = _r2_T_21 ^ _r1_T_25; // @[src/main/scala/crypto/aes/MixColumns.scala 33:34]
  wire  r2_msb_7 = bytes_15[7]; // @[src/main/scala/crypto/aes/MixColumns.scala 22:16]
  wire [8:0] _r2_sh_T_7 = {bytes_15, 1'h0}; // @[src/main/scala/crypto/aes/MixColumns.scala 23:18]
  wire [7:0] r2_sh_7 = _r2_sh_T_7[7:0]; // @[src/main/scala/crypto/aes/MixColumns.scala 23:23]
  wire [7:0] _r2_T_25 = r2_sh_7 ^ 8'h1b; // @[src/main/scala/crypto/aes/MixColumns.scala 24:17]
  wire [7:0] _r2_T_26 = r2_msb_7 ? _r2_T_25 : r2_sh_7; // @[src/main/scala/crypto/aes/MixColumns.scala 24:8]
  wire [7:0] _r2_T_27 = _r2_T_26 ^ bytes_15; // @[src/main/scala/crypto/aes/MixColumns.scala 27:38]
  wire [7:0] r2_3 = _r2_T_24 ^ _r2_T_27; // @[src/main/scala/crypto/aes/MixColumns.scala 33:45]
  wire [7:0] _r3_T_23 = _r0_T_22 ^ bytes_12; // @[src/main/scala/crypto/aes/MixColumns.scala 27:38]
  wire [7:0] _r3_T_24 = _r3_T_23 ^ bytes_13; // @[src/main/scala/crypto/aes/MixColumns.scala 34:23]
  wire [7:0] _r3_T_25 = _r3_T_24 ^ bytes_14; // @[src/main/scala/crypto/aes/MixColumns.scala 34:34]
  wire [7:0] r3_3 = _r3_T_25 ^ _r2_T_26; // @[src/main/scala/crypto/aes/MixColumns.scala 34:45]
  wire [63:0] io_out_bits_bits_lo = {r0_2,r1_2,r2_2,r3_2,r0_3,r1_3,r2_3,r3_3}; // @[src/main/scala/crypto/aes/MixColumns.scala 51:26]
  wire [63:0] io_out_bits_bits_hi = {r0,r1,r2,r3,r0_1,r1_1,r2_1,r3_1}; // @[src/main/scala/crypto/aes/MixColumns.scala 51:26]
  assign io_in_ready = io_out_ready; // @[src/main/scala/crypto/aes/MixColumns.scala 15:16]
  assign io_out_valid = io_in_valid; // @[src/main/scala/crypto/aes/MixColumns.scala 14:16]
  assign io_out_bits_bits = {io_out_bits_bits_hi,io_out_bits_bits_lo}; // @[src/main/scala/crypto/aes/MixColumns.scala 51:26]
endmodule
module AesStdRound(
  output         io_in_ready, // @[src/main/scala/crypto/aes/Round.scala 8:14]
  input          io_in_valid, // @[src/main/scala/crypto/aes/Round.scala 8:14]
  input  [127:0] io_in_bits_bits, // @[src/main/scala/crypto/aes/Round.scala 8:14]
  input  [127:0] io_rk_bits, // @[src/main/scala/crypto/aes/Round.scala 8:14]
  input          io_out_ready, // @[src/main/scala/crypto/aes/Round.scala 8:14]
  output         io_out_valid, // @[src/main/scala/crypto/aes/Round.scala 8:14]
  output [127:0] io_out_bits_bits // @[src/main/scala/crypto/aes/Round.scala 8:14]
);
  wire  sub_io_in_ready; // @[src/main/scala/crypto/aes/Round.scala 14:20]
  wire  sub_io_in_valid; // @[src/main/scala/crypto/aes/Round.scala 14:20]
  wire [127:0] sub_io_in_bits_bits; // @[src/main/scala/crypto/aes/Round.scala 14:20]
  wire  sub_io_out_ready; // @[src/main/scala/crypto/aes/Round.scala 14:20]
  wire  sub_io_out_valid; // @[src/main/scala/crypto/aes/Round.scala 14:20]
  wire [127:0] sub_io_out_bits_bits; // @[src/main/scala/crypto/aes/Round.scala 14:20]
  wire  sh_io_in_ready; // @[src/main/scala/crypto/aes/Round.scala 15:20]
  wire  sh_io_in_valid; // @[src/main/scala/crypto/aes/Round.scala 15:20]
  wire [127:0] sh_io_in_bits_bits; // @[src/main/scala/crypto/aes/Round.scala 15:20]
  wire  sh_io_out_ready; // @[src/main/scala/crypto/aes/Round.scala 15:20]
  wire  sh_io_out_valid; // @[src/main/scala/crypto/aes/Round.scala 15:20]
  wire [127:0] sh_io_out_bits_bits; // @[src/main/scala/crypto/aes/Round.scala 15:20]
  wire  mix_io_in_ready; // @[src/main/scala/crypto/aes/Round.scala 16:20]
  wire  mix_io_in_valid; // @[src/main/scala/crypto/aes/Round.scala 16:20]
  wire [127:0] mix_io_in_bits_bits; // @[src/main/scala/crypto/aes/Round.scala 16:20]
  wire  mix_io_out_ready; // @[src/main/scala/crypto/aes/Round.scala 16:20]
  wire  mix_io_out_valid; // @[src/main/scala/crypto/aes/Round.scala 16:20]
  wire [127:0] mix_io_out_bits_bits; // @[src/main/scala/crypto/aes/Round.scala 16:20]
  wire  addk_io_in_ready; // @[src/main/scala/crypto/aes/Round.scala 17:20]
  wire  addk_io_in_valid; // @[src/main/scala/crypto/aes/Round.scala 17:20]
  wire [127:0] addk_io_in_bits_bits; // @[src/main/scala/crypto/aes/Round.scala 17:20]
  wire [127:0] addk_io_rk_bits; // @[src/main/scala/crypto/aes/Round.scala 17:20]
  wire  addk_io_out_ready; // @[src/main/scala/crypto/aes/Round.scala 17:20]
  wire  addk_io_out_valid; // @[src/main/scala/crypto/aes/Round.scala 17:20]
  wire [127:0] addk_io_out_bits_bits; // @[src/main/scala/crypto/aes/Round.scala 17:20]
  SubBytes sub ( // @[src/main/scala/crypto/aes/Round.scala 14:20]
    .io_in_ready(sub_io_in_ready),
    .io_in_valid(sub_io_in_valid),
    .io_in_bits_bits(sub_io_in_bits_bits),
    .io_out_ready(sub_io_out_ready),
    .io_out_valid(sub_io_out_valid),
    .io_out_bits_bits(sub_io_out_bits_bits)
  );
  ShiftRows sh ( // @[src/main/scala/crypto/aes/Round.scala 15:20]
    .io_in_ready(sh_io_in_ready),
    .io_in_valid(sh_io_in_valid),
    .io_in_bits_bits(sh_io_in_bits_bits),
    .io_out_ready(sh_io_out_ready),
    .io_out_valid(sh_io_out_valid),
    .io_out_bits_bits(sh_io_out_bits_bits)
  );
  MixColumns mix ( // @[src/main/scala/crypto/aes/Round.scala 16:20]
    .io_in_ready(mix_io_in_ready),
    .io_in_valid(mix_io_in_valid),
    .io_in_bits_bits(mix_io_in_bits_bits),
    .io_out_ready(mix_io_out_ready),
    .io_out_valid(mix_io_out_valid),
    .io_out_bits_bits(mix_io_out_bits_bits)
  );
  AddRoundKey addk ( // @[src/main/scala/crypto/aes/Round.scala 17:20]
    .io_in_ready(addk_io_in_ready),
    .io_in_valid(addk_io_in_valid),
    .io_in_bits_bits(addk_io_in_bits_bits),
    .io_rk_bits(addk_io_rk_bits),
    .io_out_ready(addk_io_out_ready),
    .io_out_valid(addk_io_out_valid),
    .io_out_bits_bits(addk_io_out_bits_bits)
  );
  assign io_in_ready = sub_io_in_ready; // @[src/main/scala/crypto/aes/Round.scala 19:13]
  assign io_out_valid = addk_io_out_valid; // @[src/main/scala/crypto/aes/Round.scala 25:10]
  assign io_out_bits_bits = addk_io_out_bits_bits; // @[src/main/scala/crypto/aes/Round.scala 25:10]
  assign sub_io_in_valid = io_in_valid; // @[src/main/scala/crypto/aes/Round.scala 19:13]
  assign sub_io_in_bits_bits = io_in_bits_bits; // @[src/main/scala/crypto/aes/Round.scala 19:13]
  assign sub_io_out_ready = sh_io_in_ready; // @[src/main/scala/crypto/aes/Round.scala 20:13]
  assign sh_io_in_valid = sub_io_out_valid; // @[src/main/scala/crypto/aes/Round.scala 20:13]
  assign sh_io_in_bits_bits = sub_io_out_bits_bits; // @[src/main/scala/crypto/aes/Round.scala 20:13]
  assign sh_io_out_ready = mix_io_in_ready; // @[src/main/scala/crypto/aes/Round.scala 21:13]
  assign mix_io_in_valid = sh_io_out_valid; // @[src/main/scala/crypto/aes/Round.scala 21:13]
  assign mix_io_in_bits_bits = sh_io_out_bits_bits; // @[src/main/scala/crypto/aes/Round.scala 21:13]
  assign mix_io_out_ready = addk_io_in_ready; // @[src/main/scala/crypto/aes/Round.scala 22:14]
  assign addk_io_in_valid = mix_io_out_valid; // @[src/main/scala/crypto/aes/Round.scala 22:14]
  assign addk_io_in_bits_bits = mix_io_out_bits_bits; // @[src/main/scala/crypto/aes/Round.scala 22:14]
  assign addk_io_rk_bits = io_rk_bits; // @[src/main/scala/crypto/aes/Round.scala 23:14]
  assign addk_io_out_ready = io_out_ready; // @[src/main/scala/crypto/aes/Round.scala 25:10]
endmodule
module StdRoundGen(
  output         io_in_ready, // @[src/main/scala/crypto/gen/StdRoundGen.scala 13:14]
  input          io_in_valid, // @[src/main/scala/crypto/gen/StdRoundGen.scala 13:14]
  input  [127:0] io_in_bits_bits, // @[src/main/scala/crypto/gen/StdRoundGen.scala 13:14]
  input  [127:0] io_rk_bits, // @[src/main/scala/crypto/gen/StdRoundGen.scala 13:14]
  input          io_out_ready, // @[src/main/scala/crypto/gen/StdRoundGen.scala 13:14]
  output         io_out_valid, // @[src/main/scala/crypto/gen/StdRoundGen.scala 13:14]
  output [127:0] io_out_bits_bits // @[src/main/scala/crypto/gen/StdRoundGen.scala 13:14]
);
  wire  core_io_in_ready; // @[src/main/scala/crypto/gen/StdRoundGen.scala 18:20]
  wire  core_io_in_valid; // @[src/main/scala/crypto/gen/StdRoundGen.scala 18:20]
  wire [127:0] core_io_in_bits_bits; // @[src/main/scala/crypto/gen/StdRoundGen.scala 18:20]
  wire [127:0] core_io_rk_bits; // @[src/main/scala/crypto/gen/StdRoundGen.scala 18:20]
  wire  core_io_out_ready; // @[src/main/scala/crypto/gen/StdRoundGen.scala 18:20]
  wire  core_io_out_valid; // @[src/main/scala/crypto/gen/StdRoundGen.scala 18:20]
  wire [127:0] core_io_out_bits_bits; // @[src/main/scala/crypto/gen/StdRoundGen.scala 18:20]
  AesStdRound core ( // @[src/main/scala/crypto/gen/StdRoundGen.scala 18:20]
    .io_in_ready(core_io_in_ready),
    .io_in_valid(core_io_in_valid),
    .io_in_bits_bits(core_io_in_bits_bits),
    .io_rk_bits(core_io_rk_bits),
    .io_out_ready(core_io_out_ready),
    .io_out_valid(core_io_out_valid),
    .io_out_bits_bits(core_io_out_bits_bits)
  );
  assign io_in_ready = core_io_in_ready; // @[src/main/scala/crypto/gen/StdRoundGen.scala 19:14]
  assign io_out_valid = core_io_out_valid; // @[src/main/scala/crypto/gen/StdRoundGen.scala 21:10]
  assign io_out_bits_bits = core_io_out_bits_bits; // @[src/main/scala/crypto/gen/StdRoundGen.scala 21:10]
  assign core_io_in_valid = io_in_valid; // @[src/main/scala/crypto/gen/StdRoundGen.scala 19:14]
  assign core_io_in_bits_bits = io_in_bits_bits; // @[src/main/scala/crypto/gen/StdRoundGen.scala 19:14]
  assign core_io_rk_bits = io_rk_bits; // @[src/main/scala/crypto/gen/StdRoundGen.scala 20:14]
  assign core_io_out_ready = io_out_ready; // @[src/main/scala/crypto/gen/StdRoundGen.scala 21:10]
endmodule
module AesFinalRound(
  output         io_in_ready, // @[src/main/scala/crypto/aes/Round.scala 30:14]
  input          io_in_valid, // @[src/main/scala/crypto/aes/Round.scala 30:14]
  input  [127:0] io_in_bits_bits, // @[src/main/scala/crypto/aes/Round.scala 30:14]
  input  [127:0] io_rk_bits, // @[src/main/scala/crypto/aes/Round.scala 30:14]
  input          io_out_ready, // @[src/main/scala/crypto/aes/Round.scala 30:14]
  output         io_out_valid, // @[src/main/scala/crypto/aes/Round.scala 30:14]
  output [127:0] io_out_bits_bits // @[src/main/scala/crypto/aes/Round.scala 30:14]
);
  wire  sub_io_in_ready; // @[src/main/scala/crypto/aes/Round.scala 35:20]
  wire  sub_io_in_valid; // @[src/main/scala/crypto/aes/Round.scala 35:20]
  wire [127:0] sub_io_in_bits_bits; // @[src/main/scala/crypto/aes/Round.scala 35:20]
  wire  sub_io_out_ready; // @[src/main/scala/crypto/aes/Round.scala 35:20]
  wire  sub_io_out_valid; // @[src/main/scala/crypto/aes/Round.scala 35:20]
  wire [127:0] sub_io_out_bits_bits; // @[src/main/scala/crypto/aes/Round.scala 35:20]
  wire  sh_io_in_ready; // @[src/main/scala/crypto/aes/Round.scala 36:20]
  wire  sh_io_in_valid; // @[src/main/scala/crypto/aes/Round.scala 36:20]
  wire [127:0] sh_io_in_bits_bits; // @[src/main/scala/crypto/aes/Round.scala 36:20]
  wire  sh_io_out_ready; // @[src/main/scala/crypto/aes/Round.scala 36:20]
  wire  sh_io_out_valid; // @[src/main/scala/crypto/aes/Round.scala 36:20]
  wire [127:0] sh_io_out_bits_bits; // @[src/main/scala/crypto/aes/Round.scala 36:20]
  wire  addk_io_in_ready; // @[src/main/scala/crypto/aes/Round.scala 37:20]
  wire  addk_io_in_valid; // @[src/main/scala/crypto/aes/Round.scala 37:20]
  wire [127:0] addk_io_in_bits_bits; // @[src/main/scala/crypto/aes/Round.scala 37:20]
  wire [127:0] addk_io_rk_bits; // @[src/main/scala/crypto/aes/Round.scala 37:20]
  wire  addk_io_out_ready; // @[src/main/scala/crypto/aes/Round.scala 37:20]
  wire  addk_io_out_valid; // @[src/main/scala/crypto/aes/Round.scala 37:20]
  wire [127:0] addk_io_out_bits_bits; // @[src/main/scala/crypto/aes/Round.scala 37:20]
  SubBytes sub ( // @[src/main/scala/crypto/aes/Round.scala 35:20]
    .io_in_ready(sub_io_in_ready),
    .io_in_valid(sub_io_in_valid),
    .io_in_bits_bits(sub_io_in_bits_bits),
    .io_out_ready(sub_io_out_ready),
    .io_out_valid(sub_io_out_valid),
    .io_out_bits_bits(sub_io_out_bits_bits)
  );
  ShiftRows sh ( // @[src/main/scala/crypto/aes/Round.scala 36:20]
    .io_in_ready(sh_io_in_ready),
    .io_in_valid(sh_io_in_valid),
    .io_in_bits_bits(sh_io_in_bits_bits),
    .io_out_ready(sh_io_out_ready),
    .io_out_valid(sh_io_out_valid),
    .io_out_bits_bits(sh_io_out_bits_bits)
  );
  AddRoundKey addk ( // @[src/main/scala/crypto/aes/Round.scala 37:20]
    .io_in_ready(addk_io_in_ready),
    .io_in_valid(addk_io_in_valid),
    .io_in_bits_bits(addk_io_in_bits_bits),
    .io_rk_bits(addk_io_rk_bits),
    .io_out_ready(addk_io_out_ready),
    .io_out_valid(addk_io_out_valid),
    .io_out_bits_bits(addk_io_out_bits_bits)
  );
  assign io_in_ready = sub_io_in_ready; // @[src/main/scala/crypto/aes/Round.scala 38:13]
  assign io_out_valid = addk_io_out_valid; // @[src/main/scala/crypto/aes/Round.scala 42:10]
  assign io_out_bits_bits = addk_io_out_bits_bits; // @[src/main/scala/crypto/aes/Round.scala 42:10]
  assign sub_io_in_valid = io_in_valid; // @[src/main/scala/crypto/aes/Round.scala 38:13]
  assign sub_io_in_bits_bits = io_in_bits_bits; // @[src/main/scala/crypto/aes/Round.scala 38:13]
  assign sub_io_out_ready = sh_io_in_ready; // @[src/main/scala/crypto/aes/Round.scala 39:13]
  assign sh_io_in_valid = sub_io_out_valid; // @[src/main/scala/crypto/aes/Round.scala 39:13]
  assign sh_io_in_bits_bits = sub_io_out_bits_bits; // @[src/main/scala/crypto/aes/Round.scala 39:13]
  assign sh_io_out_ready = addk_io_in_ready; // @[src/main/scala/crypto/aes/Round.scala 40:14]
  assign addk_io_in_valid = sh_io_out_valid; // @[src/main/scala/crypto/aes/Round.scala 40:14]
  assign addk_io_in_bits_bits = sh_io_out_bits_bits; // @[src/main/scala/crypto/aes/Round.scala 40:14]
  assign addk_io_rk_bits = io_rk_bits; // @[src/main/scala/crypto/aes/Round.scala 41:14]
  assign addk_io_out_ready = io_out_ready; // @[src/main/scala/crypto/aes/Round.scala 42:10]
endmodule
module FinalRoundGen(
  output         io_in_ready, // @[src/main/scala/crypto/gen/FinalRoundGen.scala 13:14]
  input          io_in_valid, // @[src/main/scala/crypto/gen/FinalRoundGen.scala 13:14]
  input  [127:0] io_in_bits_bits, // @[src/main/scala/crypto/gen/FinalRoundGen.scala 13:14]
  input  [127:0] io_rk_bits, // @[src/main/scala/crypto/gen/FinalRoundGen.scala 13:14]
  input          io_out_ready, // @[src/main/scala/crypto/gen/FinalRoundGen.scala 13:14]
  output         io_out_valid, // @[src/main/scala/crypto/gen/FinalRoundGen.scala 13:14]
  output [127:0] io_out_bits_bits // @[src/main/scala/crypto/gen/FinalRoundGen.scala 13:14]
);
  wire  core_io_in_ready; // @[src/main/scala/crypto/gen/FinalRoundGen.scala 18:20]
  wire  core_io_in_valid; // @[src/main/scala/crypto/gen/FinalRoundGen.scala 18:20]
  wire [127:0] core_io_in_bits_bits; // @[src/main/scala/crypto/gen/FinalRoundGen.scala 18:20]
  wire [127:0] core_io_rk_bits; // @[src/main/scala/crypto/gen/FinalRoundGen.scala 18:20]
  wire  core_io_out_ready; // @[src/main/scala/crypto/gen/FinalRoundGen.scala 18:20]
  wire  core_io_out_valid; // @[src/main/scala/crypto/gen/FinalRoundGen.scala 18:20]
  wire [127:0] core_io_out_bits_bits; // @[src/main/scala/crypto/gen/FinalRoundGen.scala 18:20]
  AesFinalRound core ( // @[src/main/scala/crypto/gen/FinalRoundGen.scala 18:20]
    .io_in_ready(core_io_in_ready),
    .io_in_valid(core_io_in_valid),
    .io_in_bits_bits(core_io_in_bits_bits),
    .io_rk_bits(core_io_rk_bits),
    .io_out_ready(core_io_out_ready),
    .io_out_valid(core_io_out_valid),
    .io_out_bits_bits(core_io_out_bits_bits)
  );
  assign io_in_ready = core_io_in_ready; // @[src/main/scala/crypto/gen/FinalRoundGen.scala 19:14]
  assign io_out_valid = core_io_out_valid; // @[src/main/scala/crypto/gen/FinalRoundGen.scala 21:10]
  assign io_out_bits_bits = core_io_out_bits_bits; // @[src/main/scala/crypto/gen/FinalRoundGen.scala 21:10]
  assign core_io_in_valid = io_in_valid; // @[src/main/scala/crypto/gen/FinalRoundGen.scala 19:14]
  assign core_io_in_bits_bits = io_in_bits_bits; // @[src/main/scala/crypto/gen/FinalRoundGen.scala 19:14]
  assign core_io_rk_bits = io_rk_bits; // @[src/main/scala/crypto/gen/FinalRoundGen.scala 20:14]
  assign core_io_out_ready = io_out_ready; // @[src/main/scala/crypto/gen/FinalRoundGen.scala 21:10]
endmodule
module Aes128Core(
  input          clock,
  input          reset,
  output         io_in_ready, // @[src/main/scala/crypto/gen/Aes128Core.scala 18:14]
  input          io_in_valid, // @[src/main/scala/crypto/gen/Aes128Core.scala 18:14]
  input  [127:0] io_in_bits_bits, // @[src/main/scala/crypto/gen/Aes128Core.scala 18:14]
  input          io_out_ready, // @[src/main/scala/crypto/gen/Aes128Core.scala 18:14]
  output         io_out_valid, // @[src/main/scala/crypto/gen/Aes128Core.scala 18:14]
  output [127:0] io_out_bits_bits, // @[src/main/scala/crypto/gen/Aes128Core.scala 18:14]
  input  [127:0] io_key_bits // @[src/main/scala/crypto/gen/Aes128Core.scala 18:14]
);
  wire [127:0] ks_io_keyIn_bits; // @[src/main/scala/crypto/gen/Aes128Core.scala 21:18]
  wire [127:0] ks_io_rks_0_bits; // @[src/main/scala/crypto/gen/Aes128Core.scala 21:18]
  wire [127:0] ks_io_rks_1_bits; // @[src/main/scala/crypto/gen/Aes128Core.scala 21:18]
  wire [127:0] ks_io_rks_2_bits; // @[src/main/scala/crypto/gen/Aes128Core.scala 21:18]
  wire [127:0] ks_io_rks_3_bits; // @[src/main/scala/crypto/gen/Aes128Core.scala 21:18]
  wire [127:0] ks_io_rks_4_bits; // @[src/main/scala/crypto/gen/Aes128Core.scala 21:18]
  wire [127:0] ks_io_rks_5_bits; // @[src/main/scala/crypto/gen/Aes128Core.scala 21:18]
  wire [127:0] ks_io_rks_6_bits; // @[src/main/scala/crypto/gen/Aes128Core.scala 21:18]
  wire [127:0] ks_io_rks_7_bits; // @[src/main/scala/crypto/gen/Aes128Core.scala 21:18]
  wire [127:0] ks_io_rks_8_bits; // @[src/main/scala/crypto/gen/Aes128Core.scala 21:18]
  wire [127:0] ks_io_rks_9_bits; // @[src/main/scala/crypto/gen/Aes128Core.scala 21:18]
  wire [127:0] ks_io_rks_10_bits; // @[src/main/scala/crypto/gen/Aes128Core.scala 21:18]
  wire  init_io_in_ready; // @[src/main/scala/crypto/gen/Aes128Core.scala 26:20]
  wire  init_io_in_valid; // @[src/main/scala/crypto/gen/Aes128Core.scala 26:20]
  wire [127:0] init_io_in_bits_bits; // @[src/main/scala/crypto/gen/Aes128Core.scala 26:20]
  wire [127:0] init_io_rk_bits; // @[src/main/scala/crypto/gen/Aes128Core.scala 26:20]
  wire  init_io_out_ready; // @[src/main/scala/crypto/gen/Aes128Core.scala 26:20]
  wire  init_io_out_valid; // @[src/main/scala/crypto/gen/Aes128Core.scala 26:20]
  wire [127:0] init_io_out_bits_bits; // @[src/main/scala/crypto/gen/Aes128Core.scala 26:20]
  wire  r1_io_in_ready; // @[src/main/scala/crypto/gen/Aes128Core.scala 32:18]
  wire  r1_io_in_valid; // @[src/main/scala/crypto/gen/Aes128Core.scala 32:18]
  wire [127:0] r1_io_in_bits_bits; // @[src/main/scala/crypto/gen/Aes128Core.scala 32:18]
  wire [127:0] r1_io_rk_bits; // @[src/main/scala/crypto/gen/Aes128Core.scala 32:18]
  wire  r1_io_out_ready; // @[src/main/scala/crypto/gen/Aes128Core.scala 32:18]
  wire  r1_io_out_valid; // @[src/main/scala/crypto/gen/Aes128Core.scala 32:18]
  wire [127:0] r1_io_out_bits_bits; // @[src/main/scala/crypto/gen/Aes128Core.scala 32:18]
  wire  r2_io_in_ready; // @[src/main/scala/crypto/gen/Aes128Core.scala 33:18]
  wire  r2_io_in_valid; // @[src/main/scala/crypto/gen/Aes128Core.scala 33:18]
  wire [127:0] r2_io_in_bits_bits; // @[src/main/scala/crypto/gen/Aes128Core.scala 33:18]
  wire [127:0] r2_io_rk_bits; // @[src/main/scala/crypto/gen/Aes128Core.scala 33:18]
  wire  r2_io_out_ready; // @[src/main/scala/crypto/gen/Aes128Core.scala 33:18]
  wire  r2_io_out_valid; // @[src/main/scala/crypto/gen/Aes128Core.scala 33:18]
  wire [127:0] r2_io_out_bits_bits; // @[src/main/scala/crypto/gen/Aes128Core.scala 33:18]
  wire  r3_io_in_ready; // @[src/main/scala/crypto/gen/Aes128Core.scala 34:18]
  wire  r3_io_in_valid; // @[src/main/scala/crypto/gen/Aes128Core.scala 34:18]
  wire [127:0] r3_io_in_bits_bits; // @[src/main/scala/crypto/gen/Aes128Core.scala 34:18]
  wire [127:0] r3_io_rk_bits; // @[src/main/scala/crypto/gen/Aes128Core.scala 34:18]
  wire  r3_io_out_ready; // @[src/main/scala/crypto/gen/Aes128Core.scala 34:18]
  wire  r3_io_out_valid; // @[src/main/scala/crypto/gen/Aes128Core.scala 34:18]
  wire [127:0] r3_io_out_bits_bits; // @[src/main/scala/crypto/gen/Aes128Core.scala 34:18]
  wire  r4_io_in_ready; // @[src/main/scala/crypto/gen/Aes128Core.scala 35:18]
  wire  r4_io_in_valid; // @[src/main/scala/crypto/gen/Aes128Core.scala 35:18]
  wire [127:0] r4_io_in_bits_bits; // @[src/main/scala/crypto/gen/Aes128Core.scala 35:18]
  wire [127:0] r4_io_rk_bits; // @[src/main/scala/crypto/gen/Aes128Core.scala 35:18]
  wire  r4_io_out_ready; // @[src/main/scala/crypto/gen/Aes128Core.scala 35:18]
  wire  r4_io_out_valid; // @[src/main/scala/crypto/gen/Aes128Core.scala 35:18]
  wire [127:0] r4_io_out_bits_bits; // @[src/main/scala/crypto/gen/Aes128Core.scala 35:18]
  wire  r5_io_in_ready; // @[src/main/scala/crypto/gen/Aes128Core.scala 36:18]
  wire  r5_io_in_valid; // @[src/main/scala/crypto/gen/Aes128Core.scala 36:18]
  wire [127:0] r5_io_in_bits_bits; // @[src/main/scala/crypto/gen/Aes128Core.scala 36:18]
  wire [127:0] r5_io_rk_bits; // @[src/main/scala/crypto/gen/Aes128Core.scala 36:18]
  wire  r5_io_out_ready; // @[src/main/scala/crypto/gen/Aes128Core.scala 36:18]
  wire  r5_io_out_valid; // @[src/main/scala/crypto/gen/Aes128Core.scala 36:18]
  wire [127:0] r5_io_out_bits_bits; // @[src/main/scala/crypto/gen/Aes128Core.scala 36:18]
  wire  r6_io_in_ready; // @[src/main/scala/crypto/gen/Aes128Core.scala 37:18]
  wire  r6_io_in_valid; // @[src/main/scala/crypto/gen/Aes128Core.scala 37:18]
  wire [127:0] r6_io_in_bits_bits; // @[src/main/scala/crypto/gen/Aes128Core.scala 37:18]
  wire [127:0] r6_io_rk_bits; // @[src/main/scala/crypto/gen/Aes128Core.scala 37:18]
  wire  r6_io_out_ready; // @[src/main/scala/crypto/gen/Aes128Core.scala 37:18]
  wire  r6_io_out_valid; // @[src/main/scala/crypto/gen/Aes128Core.scala 37:18]
  wire [127:0] r6_io_out_bits_bits; // @[src/main/scala/crypto/gen/Aes128Core.scala 37:18]
  wire  r7_io_in_ready; // @[src/main/scala/crypto/gen/Aes128Core.scala 38:18]
  wire  r7_io_in_valid; // @[src/main/scala/crypto/gen/Aes128Core.scala 38:18]
  wire [127:0] r7_io_in_bits_bits; // @[src/main/scala/crypto/gen/Aes128Core.scala 38:18]
  wire [127:0] r7_io_rk_bits; // @[src/main/scala/crypto/gen/Aes128Core.scala 38:18]
  wire  r7_io_out_ready; // @[src/main/scala/crypto/gen/Aes128Core.scala 38:18]
  wire  r7_io_out_valid; // @[src/main/scala/crypto/gen/Aes128Core.scala 38:18]
  wire [127:0] r7_io_out_bits_bits; // @[src/main/scala/crypto/gen/Aes128Core.scala 38:18]
  wire  r8_io_in_ready; // @[src/main/scala/crypto/gen/Aes128Core.scala 39:18]
  wire  r8_io_in_valid; // @[src/main/scala/crypto/gen/Aes128Core.scala 39:18]
  wire [127:0] r8_io_in_bits_bits; // @[src/main/scala/crypto/gen/Aes128Core.scala 39:18]
  wire [127:0] r8_io_rk_bits; // @[src/main/scala/crypto/gen/Aes128Core.scala 39:18]
  wire  r8_io_out_ready; // @[src/main/scala/crypto/gen/Aes128Core.scala 39:18]
  wire  r8_io_out_valid; // @[src/main/scala/crypto/gen/Aes128Core.scala 39:18]
  wire [127:0] r8_io_out_bits_bits; // @[src/main/scala/crypto/gen/Aes128Core.scala 39:18]
  wire  r9_io_in_ready; // @[src/main/scala/crypto/gen/Aes128Core.scala 40:18]
  wire  r9_io_in_valid; // @[src/main/scala/crypto/gen/Aes128Core.scala 40:18]
  wire [127:0] r9_io_in_bits_bits; // @[src/main/scala/crypto/gen/Aes128Core.scala 40:18]
  wire [127:0] r9_io_rk_bits; // @[src/main/scala/crypto/gen/Aes128Core.scala 40:18]
  wire  r9_io_out_ready; // @[src/main/scala/crypto/gen/Aes128Core.scala 40:18]
  wire  r9_io_out_valid; // @[src/main/scala/crypto/gen/Aes128Core.scala 40:18]
  wire [127:0] r9_io_out_bits_bits; // @[src/main/scala/crypto/gen/Aes128Core.scala 40:18]
  wire  finalR_io_in_ready; // @[src/main/scala/crypto/gen/Aes128Core.scala 53:22]
  wire  finalR_io_in_valid; // @[src/main/scala/crypto/gen/Aes128Core.scala 53:22]
  wire [127:0] finalR_io_in_bits_bits; // @[src/main/scala/crypto/gen/Aes128Core.scala 53:22]
  wire [127:0] finalR_io_rk_bits; // @[src/main/scala/crypto/gen/Aes128Core.scala 53:22]
  wire  finalR_io_out_ready; // @[src/main/scala/crypto/gen/Aes128Core.scala 53:22]
  wire  finalR_io_out_valid; // @[src/main/scala/crypto/gen/Aes128Core.scala 53:22]
  wire [127:0] finalR_io_out_bits_bits; // @[src/main/scala/crypto/gen/Aes128Core.scala 53:22]
  KeySchedule ks ( // @[src/main/scala/crypto/gen/Aes128Core.scala 21:18]
    .io_keyIn_bits(ks_io_keyIn_bits),
    .io_rks_0_bits(ks_io_rks_0_bits),
    .io_rks_1_bits(ks_io_rks_1_bits),
    .io_rks_2_bits(ks_io_rks_2_bits),
    .io_rks_3_bits(ks_io_rks_3_bits),
    .io_rks_4_bits(ks_io_rks_4_bits),
    .io_rks_5_bits(ks_io_rks_5_bits),
    .io_rks_6_bits(ks_io_rks_6_bits),
    .io_rks_7_bits(ks_io_rks_7_bits),
    .io_rks_8_bits(ks_io_rks_8_bits),
    .io_rks_9_bits(ks_io_rks_9_bits),
    .io_rks_10_bits(ks_io_rks_10_bits)
  );
  AddRoundKey init ( // @[src/main/scala/crypto/gen/Aes128Core.scala 26:20]
    .io_in_ready(init_io_in_ready),
    .io_in_valid(init_io_in_valid),
    .io_in_bits_bits(init_io_in_bits_bits),
    .io_rk_bits(init_io_rk_bits),
    .io_out_ready(init_io_out_ready),
    .io_out_valid(init_io_out_valid),
    .io_out_bits_bits(init_io_out_bits_bits)
  );
  StdRoundGen r1 ( // @[src/main/scala/crypto/gen/Aes128Core.scala 32:18]
    .io_in_ready(r1_io_in_ready),
    .io_in_valid(r1_io_in_valid),
    .io_in_bits_bits(r1_io_in_bits_bits),
    .io_rk_bits(r1_io_rk_bits),
    .io_out_ready(r1_io_out_ready),
    .io_out_valid(r1_io_out_valid),
    .io_out_bits_bits(r1_io_out_bits_bits)
  );
  StdRoundGen r2 ( // @[src/main/scala/crypto/gen/Aes128Core.scala 33:18]
    .io_in_ready(r2_io_in_ready),
    .io_in_valid(r2_io_in_valid),
    .io_in_bits_bits(r2_io_in_bits_bits),
    .io_rk_bits(r2_io_rk_bits),
    .io_out_ready(r2_io_out_ready),
    .io_out_valid(r2_io_out_valid),
    .io_out_bits_bits(r2_io_out_bits_bits)
  );
  StdRoundGen r3 ( // @[src/main/scala/crypto/gen/Aes128Core.scala 34:18]
    .io_in_ready(r3_io_in_ready),
    .io_in_valid(r3_io_in_valid),
    .io_in_bits_bits(r3_io_in_bits_bits),
    .io_rk_bits(r3_io_rk_bits),
    .io_out_ready(r3_io_out_ready),
    .io_out_valid(r3_io_out_valid),
    .io_out_bits_bits(r3_io_out_bits_bits)
  );
  StdRoundGen r4 ( // @[src/main/scala/crypto/gen/Aes128Core.scala 35:18]
    .io_in_ready(r4_io_in_ready),
    .io_in_valid(r4_io_in_valid),
    .io_in_bits_bits(r4_io_in_bits_bits),
    .io_rk_bits(r4_io_rk_bits),
    .io_out_ready(r4_io_out_ready),
    .io_out_valid(r4_io_out_valid),
    .io_out_bits_bits(r4_io_out_bits_bits)
  );
  StdRoundGen r5 ( // @[src/main/scala/crypto/gen/Aes128Core.scala 36:18]
    .io_in_ready(r5_io_in_ready),
    .io_in_valid(r5_io_in_valid),
    .io_in_bits_bits(r5_io_in_bits_bits),
    .io_rk_bits(r5_io_rk_bits),
    .io_out_ready(r5_io_out_ready),
    .io_out_valid(r5_io_out_valid),
    .io_out_bits_bits(r5_io_out_bits_bits)
  );
  StdRoundGen r6 ( // @[src/main/scala/crypto/gen/Aes128Core.scala 37:18]
    .io_in_ready(r6_io_in_ready),
    .io_in_valid(r6_io_in_valid),
    .io_in_bits_bits(r6_io_in_bits_bits),
    .io_rk_bits(r6_io_rk_bits),
    .io_out_ready(r6_io_out_ready),
    .io_out_valid(r6_io_out_valid),
    .io_out_bits_bits(r6_io_out_bits_bits)
  );
  StdRoundGen r7 ( // @[src/main/scala/crypto/gen/Aes128Core.scala 38:18]
    .io_in_ready(r7_io_in_ready),
    .io_in_valid(r7_io_in_valid),
    .io_in_bits_bits(r7_io_in_bits_bits),
    .io_rk_bits(r7_io_rk_bits),
    .io_out_ready(r7_io_out_ready),
    .io_out_valid(r7_io_out_valid),
    .io_out_bits_bits(r7_io_out_bits_bits)
  );
  StdRoundGen r8 ( // @[src/main/scala/crypto/gen/Aes128Core.scala 39:18]
    .io_in_ready(r8_io_in_ready),
    .io_in_valid(r8_io_in_valid),
    .io_in_bits_bits(r8_io_in_bits_bits),
    .io_rk_bits(r8_io_rk_bits),
    .io_out_ready(r8_io_out_ready),
    .io_out_valid(r8_io_out_valid),
    .io_out_bits_bits(r8_io_out_bits_bits)
  );
  StdRoundGen r9 ( // @[src/main/scala/crypto/gen/Aes128Core.scala 40:18]
    .io_in_ready(r9_io_in_ready),
    .io_in_valid(r9_io_in_valid),
    .io_in_bits_bits(r9_io_in_bits_bits),
    .io_rk_bits(r9_io_rk_bits),
    .io_out_ready(r9_io_out_ready),
    .io_out_valid(r9_io_out_valid),
    .io_out_bits_bits(r9_io_out_bits_bits)
  );
  FinalRoundGen finalR ( // @[src/main/scala/crypto/gen/Aes128Core.scala 53:22]
    .io_in_ready(finalR_io_in_ready),
    .io_in_valid(finalR_io_in_valid),
    .io_in_bits_bits(finalR_io_in_bits_bits),
    .io_rk_bits(finalR_io_rk_bits),
    .io_out_ready(finalR_io_out_ready),
    .io_out_valid(finalR_io_out_valid),
    .io_out_bits_bits(finalR_io_out_bits_bits)
  );
  assign io_in_ready = init_io_in_ready; // @[src/main/scala/crypto/gen/Aes128Core.scala 27:14]
  assign io_out_valid = finalR_io_out_valid; // @[src/main/scala/crypto/gen/Aes128Core.scala 58:10]
  assign io_out_bits_bits = finalR_io_out_bits_bits; // @[src/main/scala/crypto/gen/Aes128Core.scala 58:10]
  assign ks_io_keyIn_bits = io_key_bits; // @[src/main/scala/crypto/gen/Aes128Core.scala 23:15]
  assign init_io_in_valid = io_in_valid; // @[src/main/scala/crypto/gen/Aes128Core.scala 27:14]
  assign init_io_in_bits_bits = io_in_bits_bits; // @[src/main/scala/crypto/gen/Aes128Core.scala 27:14]
  assign init_io_rk_bits = ks_io_rks_0_bits; // @[src/main/scala/crypto/gen/Aes128Core.scala 29:14]
  assign init_io_out_ready = r1_io_in_ready; // @[src/main/scala/crypto/gen/Aes128Core.scala 42:12]
  assign r1_io_in_valid = init_io_out_valid; // @[src/main/scala/crypto/gen/Aes128Core.scala 42:12]
  assign r1_io_in_bits_bits = init_io_out_bits_bits; // @[src/main/scala/crypto/gen/Aes128Core.scala 42:12]
  assign r1_io_rk_bits = ks_io_rks_1_bits; // @[src/main/scala/crypto/gen/Aes128Core.scala 42:37]
  assign r1_io_out_ready = r2_io_in_ready; // @[src/main/scala/crypto/gen/Aes128Core.scala 43:12]
  assign r2_io_in_valid = r1_io_out_valid; // @[src/main/scala/crypto/gen/Aes128Core.scala 43:12]
  assign r2_io_in_bits_bits = r1_io_out_bits_bits; // @[src/main/scala/crypto/gen/Aes128Core.scala 43:12]
  assign r2_io_rk_bits = ks_io_rks_2_bits; // @[src/main/scala/crypto/gen/Aes128Core.scala 43:36]
  assign r2_io_out_ready = r3_io_in_ready; // @[src/main/scala/crypto/gen/Aes128Core.scala 44:12]
  assign r3_io_in_valid = r2_io_out_valid; // @[src/main/scala/crypto/gen/Aes128Core.scala 44:12]
  assign r3_io_in_bits_bits = r2_io_out_bits_bits; // @[src/main/scala/crypto/gen/Aes128Core.scala 44:12]
  assign r3_io_rk_bits = ks_io_rks_3_bits; // @[src/main/scala/crypto/gen/Aes128Core.scala 44:36]
  assign r3_io_out_ready = r4_io_in_ready; // @[src/main/scala/crypto/gen/Aes128Core.scala 45:12]
  assign r4_io_in_valid = r3_io_out_valid; // @[src/main/scala/crypto/gen/Aes128Core.scala 45:12]
  assign r4_io_in_bits_bits = r3_io_out_bits_bits; // @[src/main/scala/crypto/gen/Aes128Core.scala 45:12]
  assign r4_io_rk_bits = ks_io_rks_4_bits; // @[src/main/scala/crypto/gen/Aes128Core.scala 45:36]
  assign r4_io_out_ready = r5_io_in_ready; // @[src/main/scala/crypto/gen/Aes128Core.scala 46:12]
  assign r5_io_in_valid = r4_io_out_valid; // @[src/main/scala/crypto/gen/Aes128Core.scala 46:12]
  assign r5_io_in_bits_bits = r4_io_out_bits_bits; // @[src/main/scala/crypto/gen/Aes128Core.scala 46:12]
  assign r5_io_rk_bits = ks_io_rks_5_bits; // @[src/main/scala/crypto/gen/Aes128Core.scala 46:36]
  assign r5_io_out_ready = r6_io_in_ready; // @[src/main/scala/crypto/gen/Aes128Core.scala 47:12]
  assign r6_io_in_valid = r5_io_out_valid; // @[src/main/scala/crypto/gen/Aes128Core.scala 47:12]
  assign r6_io_in_bits_bits = r5_io_out_bits_bits; // @[src/main/scala/crypto/gen/Aes128Core.scala 47:12]
  assign r6_io_rk_bits = ks_io_rks_6_bits; // @[src/main/scala/crypto/gen/Aes128Core.scala 47:36]
  assign r6_io_out_ready = r7_io_in_ready; // @[src/main/scala/crypto/gen/Aes128Core.scala 48:12]
  assign r7_io_in_valid = r6_io_out_valid; // @[src/main/scala/crypto/gen/Aes128Core.scala 48:12]
  assign r7_io_in_bits_bits = r6_io_out_bits_bits; // @[src/main/scala/crypto/gen/Aes128Core.scala 48:12]
  assign r7_io_rk_bits = ks_io_rks_7_bits; // @[src/main/scala/crypto/gen/Aes128Core.scala 48:36]
  assign r7_io_out_ready = r8_io_in_ready; // @[src/main/scala/crypto/gen/Aes128Core.scala 49:12]
  assign r8_io_in_valid = r7_io_out_valid; // @[src/main/scala/crypto/gen/Aes128Core.scala 49:12]
  assign r8_io_in_bits_bits = r7_io_out_bits_bits; // @[src/main/scala/crypto/gen/Aes128Core.scala 49:12]
  assign r8_io_rk_bits = ks_io_rks_8_bits; // @[src/main/scala/crypto/gen/Aes128Core.scala 49:36]
  assign r8_io_out_ready = r9_io_in_ready; // @[src/main/scala/crypto/gen/Aes128Core.scala 50:12]
  assign r9_io_in_valid = r8_io_out_valid; // @[src/main/scala/crypto/gen/Aes128Core.scala 50:12]
  assign r9_io_in_bits_bits = r8_io_out_bits_bits; // @[src/main/scala/crypto/gen/Aes128Core.scala 50:12]
  assign r9_io_rk_bits = ks_io_rks_9_bits; // @[src/main/scala/crypto/gen/Aes128Core.scala 50:36]
  assign r9_io_out_ready = finalR_io_in_ready; // @[src/main/scala/crypto/gen/Aes128Core.scala 54:16]
  assign finalR_io_in_valid = r9_io_out_valid; // @[src/main/scala/crypto/gen/Aes128Core.scala 54:16]
  assign finalR_io_in_bits_bits = r9_io_out_bits_bits; // @[src/main/scala/crypto/gen/Aes128Core.scala 54:16]
  assign finalR_io_rk_bits = ks_io_rks_10_bits; // @[src/main/scala/crypto/gen/Aes128Core.scala 55:16]
  assign finalR_io_out_ready = io_out_ready; // @[src/main/scala/crypto/gen/Aes128Core.scala 58:10]
endmodule
